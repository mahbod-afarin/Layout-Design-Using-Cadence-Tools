
module dff_0 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module and2_0 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and3_0 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and4_0 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module or2_0 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or3_0 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or4_0 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module nand2_0 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand4_0 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand3_0 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nor2_0 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor4_0 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor3_0 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module dff_1 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_2 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_3 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_4 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_5 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_6 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_7 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_8 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_9 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_10 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_11 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_12 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_13 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_14 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_15 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_16 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_17 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_18 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_19 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_20 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_21 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_22 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_23 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_24 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_25 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_26 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_27 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_28 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_29 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_30 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_31 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_32 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_33 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_34 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_35 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_36 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_37 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_38 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_39 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_40 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_41 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_42 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_43 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_44 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_45 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_46 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_47 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_48 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_49 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_50 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_51 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_52 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_53 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_54 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_55 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_56 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_57 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_58 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_59 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_60 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_61 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_62 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_63 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_64 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_65 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_66 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_67 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_68 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_69 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_70 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_71 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_72 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_73 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_74 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_75 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_76 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_77 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_78 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_79 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_80 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_81 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_82 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_83 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_84 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_85 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_86 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_87 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_88 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_89 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_90 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_91 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_92 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_93 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_94 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_95 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_96 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_97 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_98 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_99 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_100 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_101 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_102 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_103 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_104 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_105 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_106 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_107 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_108 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_109 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_110 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_111 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_112 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_113 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_114 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_115 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_116 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_117 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_118 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_119 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_120 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_121 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_122 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_123 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_124 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_125 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_126 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_127 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_128 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_129 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_130 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_131 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_132 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_133 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_134 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_135 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_136 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_137 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_138 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_139 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_140 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_141 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_142 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_143 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_144 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_145 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_146 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_147 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_148 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_149 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_150 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_151 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_152 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_153 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_154 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_155 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_156 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_157 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_158 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_159 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_160 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_161 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_162 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_163 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_164 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_165 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_166 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_167 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_168 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_169 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_170 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_171 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_172 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_173 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_174 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_175 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_176 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_177 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_178 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_179 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_180 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_181 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_182 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_183 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_184 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_185 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_186 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_187 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_188 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_189 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_190 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_191 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_192 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_193 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_194 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_195 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_196 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_197 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_198 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_199 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_200 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_201 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_202 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_203 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_204 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_205 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_206 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_207 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_208 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_209 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_210 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_211 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_212 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_213 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_214 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_215 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_216 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_217 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_218 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_219 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_220 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_221 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_222 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_223 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_224 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_225 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_226 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_227 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_228 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_229 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_230 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_231 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_232 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_233 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_234 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_235 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_236 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_237 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_238 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_239 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_240 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_241 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_242 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_243 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_244 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_245 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_246 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_247 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_248 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_249 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_250 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_251 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_252 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_253 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_254 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_255 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_256 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_257 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_258 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_259 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_260 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_261 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_262 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_263 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_264 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_265 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_266 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_267 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_268 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_269 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_270 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_271 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_272 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_273 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_274 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_275 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_276 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_277 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_278 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_279 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_280 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_281 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_282 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_283 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_284 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_285 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_286 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_287 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_288 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_289 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_290 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_291 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_292 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_293 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_294 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_295 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_296 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_297 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_298 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_299 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_300 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_301 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_302 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_303 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_304 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_305 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_306 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_307 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_308 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_309 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_310 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_311 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_312 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_313 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_314 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_315 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_316 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_317 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_318 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_319 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_320 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_321 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_322 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_323 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_324 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_325 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_326 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_327 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_328 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_329 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_330 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_331 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_332 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_333 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_334 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_335 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_336 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_337 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_338 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_339 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_340 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_341 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_342 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_343 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_344 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_345 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_346 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_347 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_348 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_349 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_350 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_351 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_352 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_353 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_354 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_355 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_356 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_357 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_358 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_359 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_360 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_361 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_362 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_363 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_364 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_365 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_366 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_367 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_368 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_369 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_370 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_371 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_372 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_373 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_374 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_375 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_376 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_377 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_378 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_379 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_380 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_381 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_382 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_383 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_384 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_385 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_386 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_387 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_388 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_389 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_390 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_391 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_392 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_393 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_394 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_395 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_396 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_397 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_398 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_399 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_400 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_401 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_402 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_403 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_404 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_405 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_406 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_407 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_408 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_409 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_410 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_411 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_412 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_413 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_414 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_415 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_416 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_417 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_418 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_419 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_420 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_421 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_422 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_423 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_424 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_425 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_426 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_427 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_428 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_429 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_430 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_431 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_432 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_433 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_434 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_435 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_436 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_437 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_438 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_439 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_440 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_441 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_442 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_443 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_444 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_445 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_446 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_447 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_448 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_449 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_450 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_451 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_452 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_453 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_454 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_455 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_456 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_457 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_458 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_459 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_460 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_461 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_462 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_463 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_464 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_465 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_466 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_467 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_468 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_469 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_470 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_471 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_472 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_473 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_474 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_475 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_476 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_477 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_478 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_479 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_480 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_481 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_482 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_483 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_484 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_485 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_486 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_487 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_488 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_489 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_490 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_491 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_492 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_493 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_494 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_495 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_496 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_497 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_498 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_499 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_500 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_501 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_502 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_503 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_504 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_505 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_506 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_507 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_508 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_509 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_510 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_511 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_512 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_513 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_514 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_515 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_516 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_517 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_518 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_519 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_520 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_521 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_522 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_523 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_524 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_525 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_526 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_527 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_528 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_529 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_530 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_531 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_532 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module dff_533 ( clk, q, d );
  input clk, d;
  output q;


  DFFHQX1 q_reg ( .D(d), .CK(clk), .Q(q) );
endmodule


module and2_1 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_2 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_3 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_4 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_5 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_6 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_7 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_8 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_9 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_10 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_11 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_12 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_13 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_14 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_15 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_16 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_17 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_18 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_19 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_20 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_21 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_22 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_23 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_24 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_25 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_26 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_27 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_28 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_29 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_30 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_31 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_32 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_33 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_34 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_35 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_36 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_37 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_38 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_39 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_40 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_41 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_42 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_43 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_44 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_45 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_46 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_47 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_48 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_49 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_50 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_51 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_52 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_53 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_54 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_55 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_56 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_57 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_58 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_59 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_60 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_61 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_62 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_63 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_64 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_65 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_66 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_67 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_68 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_69 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_70 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_71 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_72 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_73 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_74 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_75 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_76 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_77 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_78 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_79 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_80 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_81 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_82 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_83 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_84 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_85 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_86 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_87 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_88 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_89 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_90 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_91 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_92 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_93 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_94 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_95 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_96 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_97 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_98 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_99 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_100 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_101 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_102 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_103 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_104 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_105 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_106 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_107 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_108 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_109 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_110 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_111 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_112 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_113 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_114 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_115 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_116 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_117 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_118 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_119 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_120 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_121 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_122 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_123 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_124 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_125 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_126 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_127 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_128 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_129 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_130 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_131 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_132 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_133 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_134 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_135 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_136 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_137 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_138 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_139 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_140 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_141 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_142 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_143 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_144 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_145 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_146 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_147 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_148 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_149 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_150 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_151 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_152 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_153 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_154 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_155 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_156 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_157 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_158 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_159 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_160 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_161 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_162 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_163 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_164 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_165 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_166 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_167 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_168 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_169 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_170 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_171 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_172 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_173 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_174 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_175 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_176 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_177 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_178 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_179 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_180 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_181 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_182 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_183 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_184 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_185 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_186 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_187 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_188 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_189 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_190 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_191 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_192 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_193 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_194 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_195 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_196 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_197 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_198 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_199 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_200 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_201 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_202 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_203 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_204 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_205 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_206 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_207 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_208 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_209 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_210 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_211 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_212 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_213 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_214 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_215 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_216 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_217 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_218 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_219 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_220 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_221 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_222 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_223 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_224 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_225 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_226 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_227 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_228 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_229 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_230 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_231 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_232 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_233 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_234 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_235 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_236 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_237 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_238 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_239 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_240 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_241 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_242 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_243 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_244 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_245 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_246 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_247 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_248 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_249 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_250 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_251 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_252 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_253 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_254 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_255 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_256 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_257 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_258 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_259 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_260 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_261 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_262 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_263 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_264 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_265 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_266 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_267 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_268 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_269 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_270 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_271 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_272 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_273 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_274 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_275 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_276 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_277 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_278 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_279 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_280 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_281 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_282 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_283 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_284 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_285 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_286 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_287 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_288 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_289 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_290 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_291 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_292 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_293 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_294 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_295 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_296 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_297 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_298 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_299 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_300 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_301 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_302 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_303 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_304 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_305 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_306 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_307 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_308 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_309 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_310 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_311 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_312 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_313 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_314 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_315 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_316 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_317 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_318 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_319 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_320 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_321 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_322 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_323 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_324 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_325 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_326 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_327 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_328 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_329 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_330 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_331 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_332 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_333 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_334 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_335 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_336 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_337 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_338 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_339 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_340 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_341 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_342 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_343 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_344 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_345 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_346 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_347 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_348 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_349 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_350 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_351 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_352 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_353 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_354 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_355 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_356 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_357 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_358 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_359 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_360 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_361 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_362 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_363 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_364 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_365 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_366 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_367 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_368 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_369 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_370 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_371 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_372 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_373 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_374 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_375 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_376 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_377 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_378 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_379 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_380 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_381 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_382 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_383 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_384 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_385 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_386 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_387 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_388 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_389 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_390 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_391 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_392 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_393 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_394 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_395 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_396 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_397 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_398 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_399 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_400 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_401 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_402 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_403 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_404 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_405 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_406 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_407 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_408 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_409 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_410 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_411 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_412 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_413 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_414 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_415 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_416 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_417 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_418 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_419 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_420 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_421 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_422 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_423 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_424 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_425 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_426 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_427 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_428 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_429 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_430 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_431 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_432 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_433 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_434 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_435 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_436 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_437 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_438 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_439 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_440 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_441 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_442 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_443 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_444 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_445 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_446 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_447 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_448 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_449 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_450 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_451 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_452 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_453 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_454 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_455 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_456 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_457 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_458 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_459 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_460 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_461 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_462 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_463 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_464 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_465 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_466 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_467 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_468 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_469 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_470 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_471 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_472 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_473 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_474 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_475 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_476 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_477 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_478 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_479 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_480 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_481 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_482 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_483 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_484 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_485 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_486 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_487 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_488 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_489 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_490 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_491 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_492 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_493 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_494 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_495 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_496 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_497 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_498 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_499 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_500 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_501 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_502 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_503 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_504 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_505 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_506 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_507 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_508 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_509 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_510 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_511 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_512 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_513 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_514 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_515 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_516 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_517 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_518 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_519 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_520 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_521 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_522 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_523 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_524 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_525 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_526 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_527 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_528 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_529 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_530 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_531 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_532 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_533 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_534 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_535 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_536 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_537 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_538 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_539 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_540 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_541 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_542 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_543 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_544 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_545 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_546 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_547 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_548 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_549 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_550 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_551 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_552 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_553 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_554 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_555 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_556 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_557 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_558 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_559 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_560 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_561 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_562 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_563 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_564 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_565 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_566 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_567 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_568 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_569 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_570 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_571 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_572 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_573 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_574 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_575 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_576 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_577 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_578 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_579 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_580 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_581 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_582 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_583 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_584 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_585 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_586 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_587 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_588 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_589 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_590 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_591 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_592 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_593 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_594 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_595 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_596 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_597 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_598 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_599 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_600 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_601 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_602 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_603 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_604 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_605 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_606 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_607 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_608 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_609 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_610 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_611 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_612 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_613 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_614 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_615 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_616 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_617 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_618 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_619 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_620 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_621 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_622 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_623 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_624 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_625 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_626 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_627 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_628 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_629 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_630 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_631 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_632 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_633 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_634 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_635 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_636 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_637 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_638 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_639 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_640 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_641 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_642 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_643 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_644 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_645 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_646 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_647 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_648 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_649 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_650 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_651 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_652 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_653 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_654 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_655 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_656 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_657 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_658 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_659 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_660 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_661 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_662 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_663 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_664 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_665 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_666 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_667 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_668 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_669 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_670 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_671 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_672 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_673 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_674 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_675 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_676 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_677 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_678 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_679 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_680 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_681 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_682 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_683 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_684 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_685 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_686 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_687 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_688 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_689 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_690 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_691 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_692 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_693 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_694 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_695 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_696 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_697 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_698 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_699 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_700 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_701 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_702 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_703 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_704 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_705 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_706 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_707 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_708 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_709 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_710 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_711 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_712 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_713 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_714 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_715 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_716 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_717 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_718 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_719 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_720 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_721 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_722 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_723 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_724 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_725 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_726 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_727 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_728 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_729 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_730 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_731 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_732 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_733 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_734 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_735 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_736 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_737 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_738 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_739 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_740 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_741 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_742 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_743 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_744 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_745 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_746 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_747 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_748 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_749 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_750 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_751 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_752 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_753 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_754 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_755 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_756 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_757 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_758 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_759 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_760 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_761 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_762 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_763 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_764 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_765 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_766 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_767 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_768 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_769 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_770 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_771 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_772 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_773 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_774 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_775 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_776 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_777 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_778 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_779 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_780 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_781 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_782 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_783 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_784 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_785 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_786 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_787 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_788 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_789 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_790 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_791 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_792 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_793 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_794 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_795 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_796 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_797 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_798 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_799 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_800 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_801 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_802 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_803 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_804 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_805 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_806 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_807 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_808 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_809 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_810 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_811 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_812 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_813 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_814 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_815 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_816 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_817 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_818 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_819 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_820 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_821 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_822 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_823 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_824 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_825 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_826 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_827 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_828 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_829 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_830 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_831 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_832 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_833 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_834 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_835 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_836 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_837 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_838 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_839 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_840 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_841 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_842 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_843 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_844 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_845 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_846 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_847 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_848 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_849 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_850 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_851 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_852 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_853 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_854 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_855 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_856 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_857 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_858 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_859 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_860 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_861 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_862 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_863 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_864 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_865 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_866 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_867 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_868 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_869 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_870 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_871 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_872 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_873 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_874 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_875 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_876 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_877 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_878 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_879 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_880 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_881 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_882 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_883 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_884 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_885 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_886 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_887 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_888 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_889 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_890 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_891 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_892 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_893 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_894 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_895 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_896 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_897 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_898 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_899 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_900 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_901 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_902 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_903 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_904 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_905 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_906 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_907 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_908 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_909 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_910 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_911 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_912 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_913 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_914 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_915 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_916 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_917 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_918 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_919 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_920 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_921 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_922 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_923 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_924 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_925 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_926 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_927 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_928 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_929 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_930 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_931 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_932 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_933 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_934 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_935 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_936 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_937 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_938 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_939 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_940 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_941 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_942 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_943 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_944 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_945 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_946 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_947 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_948 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_949 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_950 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_951 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_952 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_953 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_954 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_955 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_956 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_957 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_958 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_959 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_960 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_961 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_962 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_963 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_964 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_965 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_966 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_967 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_968 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_969 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_970 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_971 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_972 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_973 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_974 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_975 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_976 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_977 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_978 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_979 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_980 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_981 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_982 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_983 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_984 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_985 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_986 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_987 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_988 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_989 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_990 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_991 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_992 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_993 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_994 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_995 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_996 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_997 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_998 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_999 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1000 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1001 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1002 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1003 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1004 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1005 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1006 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1007 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1008 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1009 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1010 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1011 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1012 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1013 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1014 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1015 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1016 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1017 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1018 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1019 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1020 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1021 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1022 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1023 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1024 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1025 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1026 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1027 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1028 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1029 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1030 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1031 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1032 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1033 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1034 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1035 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1036 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1037 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1038 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1039 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1040 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1041 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1042 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1043 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1044 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1045 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1046 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1047 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1048 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1049 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1050 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1051 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1052 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1053 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1054 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1055 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1056 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1057 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1058 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1059 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1060 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1061 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1062 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1063 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1064 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1065 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1066 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1067 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1068 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1069 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1070 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1071 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1072 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1073 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1074 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1075 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1076 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1077 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1078 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1079 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1080 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1081 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1082 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1083 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1084 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1085 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1086 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1087 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1088 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1089 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1090 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1091 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1092 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1093 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1094 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1095 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1096 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1097 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1098 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1099 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1100 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1101 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1102 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1103 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1104 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1105 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1106 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1107 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1108 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1109 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1110 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1111 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1112 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1113 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1114 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1115 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1116 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1117 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1118 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1119 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1120 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1121 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1122 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1123 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1124 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1125 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1126 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1127 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1128 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1129 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1130 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1131 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1132 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1133 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1134 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1135 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1136 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1137 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1138 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1139 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1140 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1141 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1142 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1143 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1144 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1145 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1146 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1147 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1148 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1149 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1150 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1151 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1152 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1153 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1154 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1155 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1156 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1157 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1158 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1159 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1160 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1161 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1162 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1163 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1164 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1165 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1166 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1167 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1168 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1169 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1170 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1171 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1172 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1173 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1174 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1175 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1176 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1177 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1178 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1179 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1180 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1181 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1182 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1183 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1184 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1185 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1186 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1187 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1188 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1189 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1190 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1191 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1192 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1193 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1194 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1195 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1196 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1197 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1198 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1199 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1200 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1201 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1202 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1203 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1204 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1205 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1206 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1207 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1208 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1209 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1210 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1211 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1212 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1213 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1214 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1215 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1216 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1217 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1218 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1219 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1220 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1221 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1222 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1223 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1224 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1225 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1226 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1227 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1228 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1229 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1230 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1231 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1232 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1233 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1234 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1235 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1236 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1237 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1238 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1239 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1240 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1241 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1242 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1243 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1244 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1245 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1246 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1247 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1248 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1249 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1250 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1251 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1252 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1253 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1254 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1255 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1256 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1257 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1258 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1259 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1260 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1261 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1262 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1263 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1264 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1265 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1266 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1267 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1268 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1269 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1270 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1271 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1272 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1273 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1274 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1275 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1276 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1277 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1278 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1279 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1280 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1281 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1282 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1283 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1284 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1285 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1286 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1287 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1288 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1289 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1290 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1291 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1292 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1293 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1294 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1295 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1296 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1297 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1298 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1299 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1300 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1301 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1302 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1303 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1304 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1305 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1306 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1307 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1308 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1309 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1310 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1311 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1312 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1313 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1314 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1315 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1316 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1317 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1318 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1319 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1320 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1321 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1322 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1323 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1324 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1325 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1326 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1327 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1328 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1329 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1330 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1331 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1332 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1333 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1334 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1335 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1336 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1337 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1338 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1339 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1340 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1341 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1342 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1343 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1344 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1345 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1346 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1347 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1348 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1349 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1350 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1351 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1352 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1353 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1354 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1355 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1356 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1357 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1358 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1359 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1360 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1361 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1362 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1363 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1364 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1365 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1366 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1367 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1368 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1369 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1370 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1371 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1372 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1373 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1374 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1375 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1376 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1377 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1378 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1379 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1380 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1381 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1382 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1383 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1384 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1385 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1386 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1387 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1388 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1389 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1390 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1391 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1392 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1393 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1394 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1395 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1396 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1397 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1398 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1399 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1400 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1401 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1402 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1403 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1404 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1405 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1406 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1407 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1408 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1409 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1410 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1411 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1412 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1413 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1414 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1415 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1416 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1417 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1418 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1419 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1420 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1421 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1422 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1423 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1424 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1425 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1426 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1427 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1428 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1429 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1430 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1431 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1432 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1433 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1434 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1435 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1436 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1437 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1438 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1439 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1440 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1441 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1442 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1443 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1444 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1445 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1446 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1447 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1448 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1449 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1450 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1451 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1452 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1453 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1454 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1455 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1456 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1457 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1458 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1459 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1460 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1461 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1462 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1463 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1464 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1465 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1466 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1467 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1468 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1469 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1470 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1471 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1472 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1473 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1474 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1475 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1476 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1477 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1478 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1479 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1480 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1481 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1482 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1483 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1484 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1485 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1486 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1487 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1488 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1489 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1490 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1491 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1492 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1493 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1494 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1495 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1496 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1497 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1498 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1499 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1500 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1501 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1502 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1503 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1504 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1505 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1506 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1507 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1508 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1509 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1510 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1511 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1512 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1513 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1514 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1515 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1516 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1517 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1518 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1519 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1520 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1521 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1522 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1523 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1524 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1525 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1526 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1527 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1528 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1529 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1530 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1531 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1532 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1533 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1534 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1535 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1536 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1537 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1538 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1539 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1540 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1541 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1542 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1543 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1544 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1545 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1546 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1547 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1548 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1549 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1550 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1551 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1552 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and2_1553 ( c, b, a );
  input b, a;
  output c;


  AND2X2 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module and3_1 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_2 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_3 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_4 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_5 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_6 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_7 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_8 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_9 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_10 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_11 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_12 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_13 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_14 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_15 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_16 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_17 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_18 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_19 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_20 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_21 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_22 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_23 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_24 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_25 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_26 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_27 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_28 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_29 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_30 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_31 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_32 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_33 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_34 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_35 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_36 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_37 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_38 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_39 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_40 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_41 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_42 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_43 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_44 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_45 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_46 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_47 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and3_48 ( d, c, b, a );
  input c, b, a;
  output d;


  AND3X2 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module and4_1 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_2 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_3 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_4 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_5 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_6 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_7 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_8 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_9 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_10 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_11 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_12 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_13 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_14 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module and4_15 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  AND4X2 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module or2_1 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_2 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_3 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_4 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_5 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_6 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_7 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_8 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_9 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_10 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_11 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_12 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_13 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_14 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_15 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_16 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_17 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_18 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_19 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_20 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_21 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_22 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_23 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_24 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_25 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_26 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_27 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_28 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_29 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_30 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_31 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_32 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_33 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_34 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_35 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_36 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_37 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_38 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_39 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_40 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_41 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_42 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_43 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_44 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_45 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_46 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_47 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_48 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_49 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_50 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_51 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_52 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_53 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_54 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_55 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_56 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_57 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_58 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_59 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_60 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_61 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_62 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_63 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_64 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_65 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_66 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_67 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_68 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_69 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_70 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_71 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_72 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_73 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_74 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_75 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_76 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_77 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_78 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_79 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_80 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_81 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_82 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_83 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_84 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_85 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_86 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_87 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_88 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_89 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_90 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_91 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_92 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_93 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_94 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_95 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_96 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_97 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_98 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_99 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_100 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_101 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_102 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_103 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_104 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_105 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_106 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_107 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_108 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_109 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_110 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_111 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_112 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_113 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_114 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_115 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_116 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_117 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_118 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_119 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_120 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_121 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_122 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_123 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_124 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_125 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_126 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_127 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_128 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_129 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_130 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_131 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_132 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_133 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_134 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_135 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_136 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_137 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_138 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_139 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_140 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_141 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_142 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_143 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_144 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_145 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_146 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_147 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_148 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_149 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_150 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_151 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_152 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_153 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_154 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_155 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_156 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_157 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_158 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_159 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_160 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_161 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_162 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_163 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_164 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_165 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_166 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_167 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_168 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_169 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_170 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_171 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_172 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_173 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_174 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_175 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_176 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_177 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_178 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_179 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_180 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_181 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_182 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_183 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_184 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_185 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_186 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_187 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_188 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_189 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_190 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_191 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_192 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_193 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_194 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_195 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_196 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_197 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_198 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_199 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_200 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_201 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_202 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_203 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_204 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_205 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_206 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_207 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_208 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_209 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_210 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_211 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_212 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_213 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_214 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_215 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_216 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_217 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_218 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_219 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_220 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_221 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_222 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_223 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_224 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_225 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_226 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_227 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_228 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_229 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_230 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_231 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_232 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_233 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_234 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_235 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_236 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_237 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_238 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_239 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_240 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_241 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_242 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_243 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_244 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_245 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_246 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_247 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_248 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_249 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_250 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_251 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_252 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_253 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_254 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_255 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_256 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_257 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_258 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_259 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_260 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_261 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_262 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_263 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_264 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_265 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_266 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_267 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_268 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_269 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_270 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_271 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_272 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_273 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_274 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_275 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_276 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_277 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_278 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_279 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_280 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_281 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_282 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_283 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_284 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_285 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_286 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_287 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_288 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_289 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_290 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_291 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_292 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_293 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_294 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_295 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_296 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_297 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_298 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_299 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_300 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_301 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_302 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_303 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_304 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_305 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_306 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_307 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_308 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_309 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_310 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_311 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_312 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_313 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_314 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_315 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_316 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_317 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_318 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_319 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_320 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_321 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_322 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_323 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_324 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_325 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_326 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_327 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_328 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_329 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_330 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_331 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_332 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_333 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_334 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_335 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_336 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_337 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_338 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_339 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_340 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_341 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_342 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_343 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_344 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_345 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_346 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_347 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_348 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_349 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_350 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_351 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_352 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_353 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_354 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_355 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_356 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_357 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_358 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_359 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_360 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_361 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_362 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_363 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_364 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_365 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_366 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_367 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_368 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_369 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_370 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_371 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_372 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_373 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_374 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_375 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_376 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_377 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_378 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_379 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_380 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_381 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_382 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_383 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_384 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_385 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_386 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_387 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_388 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_389 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_390 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_391 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_392 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_393 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_394 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_395 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_396 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_397 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_398 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_399 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_400 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_401 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_402 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_403 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_404 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_405 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_406 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_407 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_408 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_409 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_410 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_411 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_412 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_413 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_414 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_415 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_416 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_417 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_418 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_419 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_420 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_421 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_422 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_423 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_424 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_425 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_426 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_427 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_428 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_429 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_430 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_431 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_432 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_433 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_434 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_435 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_436 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_437 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_438 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_439 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_440 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_441 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_442 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_443 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_444 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_445 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_446 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_447 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_448 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_449 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_450 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_451 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_452 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_453 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_454 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_455 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_456 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_457 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_458 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_459 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_460 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_461 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_462 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_463 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_464 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_465 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_466 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_467 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_468 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_469 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_470 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_471 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_472 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_473 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_474 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_475 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_476 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_477 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_478 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_479 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_480 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_481 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_482 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_483 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_484 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_485 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_486 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_487 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_488 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_489 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_490 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_491 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_492 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_493 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_494 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_495 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_496 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_497 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_498 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_499 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_500 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_501 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_502 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_503 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_504 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_505 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_506 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_507 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_508 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_509 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_510 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_511 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_512 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_513 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_514 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_515 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_516 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_517 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_518 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_519 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_520 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_521 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_522 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_523 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_524 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_525 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_526 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_527 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_528 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_529 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_530 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_531 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_532 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_533 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_534 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_535 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_536 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_537 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_538 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_539 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_540 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_541 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_542 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_543 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_544 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_545 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_546 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_547 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_548 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_549 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_550 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_551 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_552 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_553 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_554 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_555 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_556 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_557 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_558 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_559 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_560 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_561 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_562 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_563 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_564 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_565 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_566 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_567 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_568 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_569 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_570 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_571 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_572 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_573 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_574 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_575 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_576 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_577 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_578 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_579 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_580 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_581 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_582 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_583 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_584 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_585 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or2_586 ( c, b, a );
  input b, a;
  output c;


  OR2X2 U1 ( .A(a), .B(b), .Y(c) );
endmodule


module or3_1 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_2 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_3 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_4 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_5 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_6 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_7 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_8 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_9 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_10 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_11 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_12 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_13 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_14 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_15 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_16 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_17 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_18 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_19 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_20 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_21 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_22 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_23 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_24 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_25 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_26 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_27 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_28 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_29 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_30 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_31 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_32 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_33 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_34 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_35 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_36 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_37 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_38 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_39 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_40 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_41 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_42 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_43 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_44 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_45 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_46 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_47 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_48 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_49 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_50 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_51 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_52 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_53 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_54 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_55 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_56 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_57 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_58 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_59 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_60 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or3_61 ( d, c, b, a );
  input c, b, a;
  output d;


  OR3XL U1 ( .A(c), .B(b), .C(a), .Y(d) );
endmodule


module or4_1 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_2 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_3 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_4 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_5 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_6 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_7 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_8 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_9 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_10 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_11 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_12 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_13 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_14 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_15 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_16 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_17 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_18 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_19 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_20 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_21 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_22 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_23 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_24 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_25 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_26 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_27 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_28 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_29 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_30 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_31 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_32 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_33 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_34 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_35 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_36 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_37 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_38 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_39 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_40 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_41 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_42 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_43 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_44 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_45 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_46 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_47 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_48 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_49 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_50 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_51 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_52 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_53 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_54 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_55 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_56 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_57 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_58 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_59 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module or4_60 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  OR4X2 U1 ( .A(b), .B(a), .C(d), .D(c), .Y(e) );
endmodule


module nand2_1 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_2 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_3 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_4 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_5 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_6 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_7 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_8 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_9 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_10 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_11 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_12 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_13 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_14 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_15 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_16 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_17 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_18 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_19 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_20 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_21 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_22 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_23 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_24 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_25 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_26 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_27 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_28 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_29 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_30 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_31 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_32 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_33 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_34 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_35 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_36 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_37 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_38 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_39 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_40 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_41 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_42 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_43 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_44 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_45 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_46 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_47 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_48 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_49 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_50 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_51 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_52 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_53 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_54 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_55 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_56 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_57 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_58 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_59 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_60 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_61 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_62 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_63 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_64 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_65 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_66 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_67 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_68 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_69 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_70 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_71 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_72 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_73 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_74 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_75 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_76 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_77 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_78 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_79 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_80 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_81 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_82 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_83 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_84 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_85 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_86 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_87 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_88 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_89 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_90 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_91 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_92 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_93 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_94 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_95 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_96 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_97 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_98 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_99 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_100 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_101 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_102 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_103 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_104 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_105 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_106 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_107 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_108 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_109 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_110 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_111 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_112 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_113 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_114 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_115 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_116 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_117 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_118 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_119 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_120 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_121 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_122 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_123 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_124 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_125 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_126 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_127 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_128 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_129 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_130 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_131 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_132 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_133 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_134 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_135 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_136 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_137 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_138 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_139 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_140 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_141 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_142 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_143 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_144 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_145 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_146 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_147 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_148 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_149 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_150 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_151 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_152 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_153 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_154 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_155 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_156 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_157 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_158 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_159 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_160 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_161 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_162 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_163 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_164 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_165 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_166 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_167 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_168 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_169 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_170 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_171 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_172 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_173 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_174 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_175 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_176 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_177 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_178 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_179 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_180 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_181 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_182 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_183 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_184 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_185 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_186 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_187 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_188 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_189 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_190 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_191 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_192 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_193 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_194 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_195 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_196 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_197 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_198 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_199 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_200 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_201 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_202 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_203 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_204 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_205 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_206 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_207 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_208 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_209 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_210 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_211 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_212 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_213 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_214 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_215 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_216 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_217 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_218 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_219 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_220 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_221 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_222 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_223 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_224 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_225 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_226 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_227 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_228 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_229 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_230 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_231 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_232 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_233 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_234 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_235 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_236 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_237 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_238 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_239 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_240 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_241 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_242 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_243 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_244 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_245 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_246 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_247 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_248 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_249 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_250 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_251 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_252 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_253 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_254 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_255 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_256 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_257 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_258 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_259 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_260 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_261 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_262 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_263 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_264 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_265 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_266 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_267 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_268 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_269 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_270 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_271 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_272 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_273 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_274 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_275 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_276 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_277 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_278 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_279 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_280 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_281 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_282 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_283 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_284 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_285 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_286 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_287 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_288 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_289 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_290 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_291 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_292 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_293 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_294 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_295 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_296 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_297 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_298 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_299 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_300 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_301 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_302 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_303 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_304 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_305 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_306 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_307 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_308 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_309 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_310 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_311 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_312 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_313 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_314 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_315 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_316 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_317 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_318 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_319 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_320 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_321 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_322 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_323 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_324 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_325 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_326 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_327 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_328 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_329 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_330 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_331 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_332 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_333 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_334 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_335 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_336 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_337 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_338 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_339 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_340 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_341 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_342 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_343 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_344 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_345 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_346 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_347 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_348 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_349 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_350 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_351 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_352 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_353 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_354 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_355 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_356 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_357 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_358 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_359 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_360 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_361 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_362 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_363 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_364 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_365 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_366 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_367 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_368 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_369 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_370 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_371 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_372 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_373 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_374 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_375 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_376 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_377 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_378 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_379 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_380 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_381 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_382 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_383 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_384 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_385 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_386 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_387 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_388 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_389 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_390 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_391 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_392 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_393 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_394 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_395 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_396 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_397 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_398 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_399 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_400 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_401 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_402 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_403 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_404 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_405 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_406 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_407 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_408 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_409 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_410 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_411 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_412 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_413 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_414 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_415 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_416 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_417 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_418 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_419 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_420 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_421 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_422 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_423 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_424 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_425 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_426 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_427 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_428 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_429 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_430 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_431 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_432 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_433 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_434 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_435 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_436 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_437 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_438 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_439 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_440 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_441 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_442 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_443 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_444 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_445 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_446 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_447 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_448 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_449 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_450 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_451 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_452 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_453 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_454 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_455 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_456 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_457 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_458 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_459 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_460 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_461 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_462 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_463 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_464 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_465 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_466 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_467 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_468 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_469 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_470 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_471 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_472 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_473 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_474 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_475 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_476 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_477 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_478 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_479 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_480 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_481 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_482 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_483 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_484 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_485 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_486 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_487 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_488 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_489 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_490 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_491 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_492 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_493 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_494 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_495 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_496 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_497 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_498 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_499 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_500 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_501 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_502 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_503 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_504 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_505 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_506 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_507 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_508 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_509 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_510 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_511 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_512 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_513 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_514 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_515 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_516 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_517 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_518 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_519 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_520 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_521 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_522 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_523 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_524 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_525 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_526 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_527 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_528 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_529 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_530 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_531 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_532 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_533 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_534 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_535 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_536 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_537 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_538 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_539 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_540 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_541 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_542 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_543 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_544 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_545 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_546 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_547 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_548 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_549 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_550 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_551 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_552 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_553 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_554 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_555 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_556 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_557 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_558 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_559 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_560 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_561 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_562 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_563 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_564 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_565 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_566 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_567 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_568 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_569 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_570 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_571 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_572 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_573 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_574 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_575 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_576 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_577 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_578 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_579 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_580 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_581 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_582 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_583 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_584 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_585 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_586 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_587 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_588 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_589 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_590 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_591 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_592 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_593 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_594 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_595 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_596 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_597 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_598 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_599 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_600 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_601 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_602 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_603 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_604 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_605 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_606 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_607 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_608 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_609 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_610 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_611 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_612 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_613 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_614 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_615 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_616 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_617 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_618 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_619 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_620 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_621 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_622 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_623 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_624 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_625 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_626 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_627 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_628 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_629 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_630 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_631 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_632 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_633 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_634 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_635 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_636 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_637 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_638 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_639 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_640 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_641 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_642 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_643 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_644 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_645 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_646 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_647 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_648 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_649 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_650 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_651 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_652 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_653 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_654 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_655 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_656 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_657 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_658 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_659 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_660 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_661 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_662 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_663 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_664 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_665 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_666 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_667 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_668 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_669 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_670 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_671 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_672 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_673 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_674 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_675 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_676 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_677 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_678 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_679 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_680 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_681 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_682 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_683 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_684 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_685 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_686 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_687 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_688 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_689 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_690 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_691 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_692 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_693 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_694 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_695 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_696 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_697 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_698 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_699 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_700 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_701 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_702 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_703 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_704 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_705 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_706 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_707 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_708 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_709 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_710 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_711 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_712 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_713 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_714 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_715 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_716 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_717 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_718 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_719 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_720 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_721 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_722 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_723 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_724 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_725 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_726 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_727 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_728 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_729 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_730 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_731 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_732 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_733 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_734 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_735 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_736 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_737 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_738 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_739 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_740 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_741 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_742 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_743 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_744 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_745 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_746 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_747 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_748 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_749 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_750 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_751 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_752 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_753 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_754 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_755 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_756 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_757 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_758 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_759 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_760 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_761 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_762 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_763 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_764 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_765 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_766 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_767 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_768 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_769 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_770 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_771 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_772 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_773 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_774 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_775 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_776 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_777 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_778 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_779 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_780 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_781 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_782 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_783 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_784 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_785 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_786 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_787 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_788 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_789 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_790 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_791 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_792 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_793 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_794 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_795 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_796 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_797 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_798 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_799 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_800 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_801 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_802 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_803 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_804 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_805 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_806 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_807 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_808 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_809 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_810 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_811 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_812 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_813 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_814 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_815 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_816 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_817 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_818 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_819 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_820 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_821 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_822 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_823 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_824 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_825 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_826 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_827 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_828 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_829 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_830 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_831 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_832 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_833 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_834 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_835 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_836 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_837 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_838 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_839 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_840 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_841 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_842 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_843 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_844 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_845 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_846 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_847 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_848 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_849 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_850 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_851 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_852 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_853 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_854 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_855 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_856 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_857 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_858 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_859 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_860 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_861 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_862 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_863 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_864 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_865 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_866 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_867 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_868 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_869 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_870 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_871 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_872 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_873 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_874 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_875 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_876 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_877 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_878 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_879 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_880 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_881 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_882 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_883 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_884 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_885 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_886 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_887 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_888 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_889 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_890 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_891 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_892 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_893 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_894 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_895 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_896 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_897 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_898 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_899 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_900 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_901 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_902 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_903 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_904 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_905 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_906 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_907 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_908 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_909 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_910 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_911 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_912 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_913 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_914 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_915 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_916 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_917 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_918 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_919 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_920 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_921 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_922 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand2_923 ( c, b, a );
  input b, a;
  output c;


  NAND2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nand4_1 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_2 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_3 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_4 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_5 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_6 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_7 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_8 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_9 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_10 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_11 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_12 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_13 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_14 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_15 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_16 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_17 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_18 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_19 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand4_20 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NAND4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nand3_1 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_2 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_3 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_4 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_5 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_6 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_7 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_8 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_9 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_10 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_11 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_12 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_13 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_14 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_15 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_16 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_17 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_18 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_19 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_20 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_21 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nand3_22 ( d, c, b, a );
  input c, b, a;
  output d;


  NAND3X1 U1 ( .A(b), .B(a), .C(c), .Y(d) );
endmodule


module nor2_1 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_2 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_3 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_4 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_5 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_6 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_7 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_8 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_9 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_10 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_11 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_12 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_13 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_14 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_15 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_16 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_17 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_18 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_19 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_20 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_21 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_22 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_23 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_24 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_25 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_26 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_27 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_28 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_29 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_30 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_31 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_32 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_33 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_34 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_35 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_36 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_37 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_38 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_39 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_40 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_41 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_42 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_43 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_44 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_45 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_46 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_47 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_48 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_49 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_50 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_51 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_52 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_53 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_54 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_55 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_56 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_57 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_58 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_59 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_60 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_61 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_62 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_63 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_64 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_65 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_66 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_67 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_68 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_69 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_70 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_71 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_72 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_73 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_74 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_75 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_76 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_77 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_78 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_79 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_80 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_81 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_82 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_83 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_84 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_85 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_86 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_87 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_88 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_89 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_90 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_91 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_92 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_93 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_94 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_95 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_96 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor2_97 ( c, b, a );
  input b, a;
  output c;


  NOR2X1 U1 ( .A(b), .B(a), .Y(c) );
endmodule


module nor4_1 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_2 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_3 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_4 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_5 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_6 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_7 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_8 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_9 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_10 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_11 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_12 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_13 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_14 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_15 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_16 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_17 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_18 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_19 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_20 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_21 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_22 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_23 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_24 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_25 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_26 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_27 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_28 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_29 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_30 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_31 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_32 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_33 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_34 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_35 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_36 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_37 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_38 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_39 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_40 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor4_41 ( e, d, c, b, a );
  input d, c, b, a;
  output e;


  NOR4X1 U1 ( .A(d), .B(c), .C(b), .D(a), .Y(e) );
endmodule


module nor3_1 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_2 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_3 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_4 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_5 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_6 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_7 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_8 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_9 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module nor3_10 ( d, c, b, a );
  input c, b, a;
  output d;


  NOR3X1 U1 ( .A(a), .B(c), .C(b), .Y(d) );
endmodule


module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1960, g1961, g27,
         g28, g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g82, g83,
         g84, g85, g86, g87, g872, g873, g88, g886, g889, g89, g892, g895,
         g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92, g922,
         g925, g93, g94, g95, g96, g99, g1289, g1882, g312, g452, g11257, g123,
         g207, g713, g1153, g1209, g1744, g1558, g695, g461, g940, g976, g709,
         g8432, g1092, g1574, g1864, g369, g1580, g1736, g39, g1651, g1424,
         g1737, g1672, g1077, g1231, g4, g774, g1104, g1304, g7290, g243,
         g1499, g1044, g1444, g757, g786, g1543, g552, g315, g1534, g622,
         g1927, g1660, g278, g1436, g718, g8433, g76, g554, g496, g11333, g981,
         g878, g590, g829, g1095, g704, g1265, g7302, g1786, g682, g8429,
         g1296, g7292, g587, g52, g646, g327, g1389, g1371, g1956, g1955,
         g1675, g354, g113, g639, g1684, g1639, g1791, g248, g1707, g1759,
         g351, g1604, g1098, g932, g126, g1896, g8282, g736, g8435, g1019,
         g1362, g745, g1419, g58, g32, g876, g1086, g1486, g1730, g1504, g1470,
         g822, g583, g1678, g174, g1766, g1801, g186, g959, g1169, g1007,
         g1407, g1059, g1868, g758, g1718, g396, g11265, g1015, g38, g632,
         g1415, g1227, g1721, g882, g883, g16, g284, g426, g11256, g219, g1216,
         g1360, g806, g1428, g579, g1564, g1741, g225, g281, g1308, g611, g631,
         g1217, g1589, g1466, g1571, g1861, g1365, g1448, g1711, g1133, g1333,
         g153, g962, g766, g588, g486, g11331, g471, g1397, g580, g1950, g8288,
         g756, g755, g635, g1101, g549, g1041, g105, g1669, g1368, g1531,
         g1458, g572, g1011, g33, g1411, g1074, g444, g11259, g1474, g1080,
         g1713, g333, g269, g401, g11266, g1857, g9, g664, g965, g1400, g309,
         g814, g231, g557, g586, g869, g875, g1383, g158, g627, g1023, g259,
         g1361, g1206, g1327, g654, g293, g1346, g1633, g1753, g1508, g1240,
         g7297, g538, g11326, g416, g11269, g542, g11325, g1681, g374, g563,
         g1914, g8284, g530, g11328, g575, g1936, g55, g1117, g1317, g1356,
         g357, g386, g11263, g1601, g553, g166, g501, g11334, g262, g1840, g70,
         g318, g794, g36, g302, g342, g1250, g7299, g1163, g1810, g1032, g1432,
         g1053, g1453, g363, g330, g1157, g1357, g35, g928, g261, g516, g11337,
         g254, g778, g861, g1627, g1292, g7293, g290, g1850, g770, g1583, g466,
         g1561, g1527, g1546, g287, g560, g617, g17, g336, g456, g305, g345,
         g8, g1771, g865, g255, g1945, g1738, g1478, g1035, g1959, g1690,
         g1482, g1110, g296, g1663, g700, g8431, g1762, g360, g192, g1657,
         g722, g61, g566, g1394, g1089, g1071, g986, g971, g143, g1814, g1038,
         g1212, g1918, g782, g1822, g237, g746, g1062, g1462, g178, g366, g837,
         g599, g1854, g944, g1941, g8287, g170, g1520, g686, g953, g1958, g40,
         g1765, g1733, g1270, g7303, g1610, g1796, g1324, g1540, g1377, g491,
         g11332, g1849, g213, g1781, g1900, g1245, g7298, g108, g630, g148,
         g833, g1923, g8285, g936, g1215, g1314, g849, g1336, g272, g1806,
         g826, g1065, g1887, g8281, g37, g968, g1845, g1137, g1891, g1255,
         g7300, g257, g874, g591, g731, g636, g1218, g605, g79, g182, g950,
         g1129, g857, g448, g11258, g1828, g1727, g1592, g1703, g1932, g8286,
         g1624, g26, g1068, g578, g440, g11260, g476, g11338, g119, g668, g139,
         g1149, g34, g1848, g263, g818, g1747, g802, g275, g1524, g1577, g810,
         g391, g11264, g658, g1386, g253, g1125, g201, g1280, g7295, g1083,
         g650, g1636, g853, g421, g11270, g762, g956, g378, g1756, g589, g841,
         g1027, g1003, g1403, g1145, g1107, g1223, g406, g11267, g1811, g1642,
         g1047, g1654, g197, g1595, g1537, g727, g8434, g999, g798, g481,
         g11324, g754, g1330, g845, g790, g1512, g114, g1490, g1166, g1056,
         g348, g868, g1260, g7301, g260, g131, g7, g258, g521, g11330, g1318,
         g1872, g677, g582, g1393, g1549, g947, g1834, g1598, g1121, g1321,
         g506, g11335, g546, g1909, g1552, g584, g1687, g1586, g324, g1141,
         g1570, g1341, g1710, g1645, g115, g135, g525, g11329, g581, g1607,
         g321, g67, g1275, g11443, g1311, g1615, g382, g1374, g266, g1284,
         g7294, g1380, g673, g8428, g1853, g162, g411, g11268, g431, g11262,
         g1905, g8283, g1515, g1630, g49, g991, g1300, g7291, g339, g256,
         g1750, g585, g1440, g1666, g1528, g1351, g1648, g127, g1618, g1235,
         g7296, g299, g435, g11261, g64, g1555, g995, g1621, g1113, g643,
         g1494, g1567, g691, g8430, g534, g11327, g1776, g569, g1160, g1050,
         g1, g511, g11336, g1724, g12, g1878, g73, g4500, g5529, g9968, g4682,
         g2807, g4130, g5024, g4338, g8147, g6551, g10865, g8054, g9974, g7709,
         g4940, g4640, g4565, g11519, g5935, g4736, g6481, g6215, g10563,
         g5013, g11221, g5212, g6529, g5008, g3829, g9995, g10707, g3435,
         g5576, g10013, g10385, g3753, g4722, g9696, g10408, g10937, g7242,
         g10336, g5229, g8940, g4560, g10855, g7996, g3586, g10496, g3399,
         g6907, g8226, g5405, g6155, g7246, g6638, g11647, g2744, g3374, g8814,
         g10950, g5477, g6910, g10417, g6488, g7712, g6828, g7638, g3015,
         g10800, g4300, g8019, g6821, g8267, g11478, g3698, g4144, g3992,
         g4585, g7934, g6516, g8244, g4753, g8631, g4807, g10793, g5910, g9454,
         g2563, g2478, g3215, g10726, g6824, g9931, g5361, g10558, g5248,
         g3880, g5557, g6759, g6502, g10797, g8241, g4471, g10780, g11625,
         g11372, g10007, g10771, g9720, g5803, g11231, g11580, g5478, g4998,
         g10019, g4114, g11293, g4779, g5820, g8173, g3111, g4977, g6533,
         g3688, g5867, g10405, g7932, g10448, g5001, g8245, g8451, g8214,
         g3041, g10767, g10599, g10501, g8512, g2276, g6000, g10809, g11492,
         g4490, g8488, g4903, g10720, g10334, g6934, g5309, g6123, g6838,
         g4905, g10798, g10785, g8187, g7204, g6830, g8944, g5543, g5300,
         g8921, g8745, g6096, g6003, g3431, g10740, g6733, g6548, g5502, g6823,
         g4890, g3381, g10863, g8039, g6526, g10664, g7189, g5278, g8923,
         g5173, g10712, g4264, g6755, g2791, g5226, g11514, g10411, g4506,
         g10348, g9324, g10001, g5526, g4788, g4465, g8289, g8203, g5403,
         g6902, g6015, g11340, g6542, g4537, g6507, g10485, g5556, g8505,
         g8603, g11641, g3423, g10765, g4801, g11305, g6126, g5493, g10414,
         g7986, g8000, g10522, g8060, g7191, g8746, g10557, g5150, g6469,
         g10452, g4498, g8744, g5514, g6627, g4893, g10268, g9257, g5194,
         g3418, g6901, g8043, g5263, g6929, g5857, g8049, g4529, g9699, g6786,
         g7218, g6234, g5824, g7101, g10864, g7651, g8816, g10862, g11077,
         g3222, g3101, g9268, g5942, g10331, g10721, g8051, g10383, g6541,
         g9088, g10773, g8193, g6523, g8546, g5404, g11393, g5258, g8265,
         g2984, g11561, g4765, g4334, g11233, g7950, g6908, g8768, g8885,
         g5271, g6333, g10515, g6045, g7590, g6468, g10782, g10886, g6672,
         g6840, g5230, g8743, g3354, g5914, g7705, g7953, g10025, g6038, g4488,
         g3863, g6471, g11303, g5266, g10663, g8920, g4283, g10788, g4484,
         g8815, g3008, g9713, g4770, g5842, g7671, g5396, g7203, g10382,
         g10583, g8045, g7843, g8269, g3104, g3425, g6537, g5221, g4902, g6080,
         g5485, g6059, g4089, g7664, g8551, g5126, g10866, g10597, g11603,
         g6332, g4231, g11249, g10779, g11488, g3438, g5354, g5295, g5918,
         g6894, g3513, g4076, g6534, g6928, g3414, g8055, g11291, g3209, g6833,
         g6918, g6915, g6911, g8812, g4553, g7441, g5996, g8047, g6653, g6832,
         g4771, g11481, g10857, g7947, g3681, g6478, g4117, g6897, g6042,
         g11229, g10402, g4342, g4330, g8221, g11609, g10859, g6054, g6508,
         g6531, g8050, g8261, g11376, g8559, g2260, g10556, g7032, g8390,
         g4548, g4293, g5390, g4561, g8200, g8767, g3071, g7987, g4480, g11483,
         g10702, g5863, g5392, g5838, g8270, g10776, g6513, g9272, g10732,
         g10898, g8052, g4325, g4421, g5319, g8766, g10555, g6205, g8820,
         g9124, g6839, g6522, g10936, g11320, g6841, g10328, g8769, g6224,
         g11349, g6470, g11225, g5755, g6515, g3003, g9710, g3631, g5182,
         g11430, g10791, g5004, g7632, g11485, g6331, g5257, g8053, g4518,
         g4764, g5763, g6480, g6795, g8194, g2257, g5201, g5269, g8938, g7990,
         g4238, g8775, g4891, g8266, g11290, g6501, g10570, g6334, g10719,
         g4727, g4274, g8765, g6916, g8811, g5174, g11308, g5847, g10554,
         g10784, g2979, g10396, g11425, g7062, g5548, g6820, g4340, g6922,
         g6747, g11391, g8818, g8649, g9555, g6071, g7942, g10858, g8926,
         g4239, g11602, g8041, g8922, g5536, g5810, g7067, g8236, g11605,
         g8048, g6528, g6524, g3056, g7258, g7219, g8046, g3706, g11482,
         g10381, g4477, g10333, g2310, g6923, g4255, g4732, g8937, g4752,
         g6538, g10339, g3524, g11306, g7183, g4778, g6895, g11223, g6163,
         g6179, g9052, g9721, g8776, g6827, g4309, g9331, g7244, g7586, g7930,
         g11300, g10718, g5445, g11227, g6088, g8206, g6679, g11636, g11219,
         g2117, g3062, g9266, g11608, g8059, g8771, g2459, g6035, g7106, g6198,
         g7992, g8973, g6834, g5148, g7134, g10795, g11276, g10770, g9271,
         g10494, g8773, g3462, g3662, g6740, g10484, g7143, g8939, g8772,
         g6093, g6500, g10500, g2794, g6485, g8777, g6244, g5304, g11640,
         g4784, g11487, g9110, g11380, g9269, g7054, g7236, g3247, g11314,
         g5276, g9150, g11298, g7202, g6819, g2987, g5317, g10453, g6243,
         g6514, g8817, g8810, g9313, g6983, g8366, g4473, g6577, g3200, g8040,
         g5255, g6900, g8042, g11490, g8230, g6546, g8574, g5770, g8889,
         g10711, g9719, g11312, g5287, g6351, g6479, g3120, g5814, g5849,
         g10559, g5219, g7240, g8819, g9256, g6656, g6906, g10717, g4759,
         g5189, g8770, g6392, g6621, g11610, g4582, g8264, g11604, g2161,
         g7245, g2510, g2439, g11486, g7581, g10799, g10357, g6439, g8507,
         g7133, g8642, g8044, g8254, g11549, g11232, g11607, g6573, g3506,
         g3407, g6193, g3108, g7225, g7231, g4576, g4904, g8806, g11292, g6822,
         g7624, g3661, g6912, g6898, g5421, g7994, g8813, g6924, g5308, g11310,
         g11294, g5852, g2970, g6026, g10369, g5286, g4554, g8024, g8945,
         g4804, g6525, g6019, g8210, g5083, g3585, g7541, g4760, g10860,
         g10502, g11579, g11639, g5030, g6826, g2303, g7626, g6829, g7211,
         g7660, g10722, g8887, g11484, g11286, g6002, g11606, g11217, g10454,
         g6757, g6216, g8941, g10856, g4892, g6930, g8250, g5250, g6049, g8943,
         g10861, g8779, g5484, g3304, g4482, g5190, g6180, g5274, g8774,
         g10325, g8260, g6099, g10401, g6831, g6068, g7137, g6545, g7257,
         g6909, g8384, g11392, g6506, g8883, g6728, g10724, g4556, g3070,
         g11103, g2250, g9900, g11095, g4973, g7389, g7888, g7465, g4969,
         g8224, g2892, g5686, g10308, g4123, g8120, g6788, g5598, g4824, g9694,
         g10495, g2945, g11190, g8789, g8639, g9852, g9728, g9563, g5625,
         g4875, g9701, g7138, g10752, g11211, g11058, g11024, g8547, g8307,
         g10669, g7707, g4884, g3813, g4839, g9870, g6640, g9650, g9240, g5687,
         g7957, g3512, g7449, g4235, g4343, g11296, g9594, g9292, g9943, g9923,
         g9367, g5525, g8876, g10705, g10564, g9934, g9913, g9624, g6225,
         g6324, g10686, g6540, g8663, g11581, g6206, g3989, g7730, g7260,
         g7504, g7185, I5689, I5690, g7881, g11070, g9859, g9736, g9573, g8877,
         g11590, g2274, g6199, g8932, g5545, g5180, g5591, g8556, g8412,
         g11094, g5853, g5044, g6245, g4360, g8930, g5507, g11150, g3087,
         g8464, g8302, g9692, g4996, g7131, g11019, g9960, g9951, g9536,
         g11196, g11018, g10595, g10550, g10433, g10623, g10544, g4878, g5204,
         g4838, g8844, g8609, g6701, g6185, g10725, g5100, g4882, g8731, g5128,
         g6886, g8557, g8415, g8966, g8071, g11597, g9828, g9722, g9785, g2918,
         g9830, g9725, g8955, g9592, g5123, g7059, g6078, g7459, g11102, g7718,
         g7535, g9703, g5528, g5151, g9932, g9911, g5530, g2760, g8629, g6887,
         g6187, g6228, g5605, g6322, I6337, I6338, g8967, g5010, g3275, g2895,
         g7721, g9866, g9716, g10808, g10744, g3047, g4492, g3685, g8822,
         g8614, g10560, g11456, g9848, g9724, g9557, g4714, g6550, g5172,
         g10642, g3284, g2531, g9855, g5618, g6891, g7940, g11085, g4968,
         g8837, g8646, g9644, g9125, g5804, g8462, g8300, I6330, g11156, g6342,
         g9867, g9717, g4871, g10435, g7741, g9386, g9151, g8842, g8607, g9599,
         g9274, g8974, g5518, g9614, g9111, g4122, g7217, g4610, g11557, g2911,
         g11210, g7466, g9939, g9918, g11279, g10518, g10513, g10440, I16145,
         g8708, g7055, g5264, g6329, g8176, g8005, g7510, g4099, g3281, g11601,
         g11187, g6746, g6221, g8630, g9622, g11143, g10923, g9904, g9886,
         g9676, g8733, g6624, g11169, g8073, g9841, g9706, g9512, g5882, g5592,
         g8796, g8645, g11168, g4269, g5611, g8069, g9695, g10304, g8469,
         g8305, g4712, g6576, g5762, g10622, g11015, g5217, g5674, g9359,
         g9173, g9223, g8960, g11556, g9858, g5541, g4534, g5897, g6699, g6177,
         g6855, g3804, g3098, g5680, g9642, g5744, g8399, g9447, g9030, g11178,
         g8510, g8414, g6319, g11186, g3908, g2951, g6352, g9595, g9205, g4831,
         g4109, g5492, g8934, g10312, g6186, g9612, g9417, g9935, g9914, g8701,
         g10745, g10658, g11216, g9328, g8971, g11587, g6325, g7368, g6083,
         g6544, g5476, g7743, g4869, g5722, g6790, g5813, g8408, g10761, g7734,
         g8136, g7926, g5569, g9902, g9392, g8623, g5500, g2496, g6756, g3010,
         g5877, g8972, g6622, g11612, g9366, g11230, g4364, g9649, g5795,
         g5737, g4054, g6345, g5823, g11275, g9851, g6763, g5802, I16142,
         g10511, g10509, g10507, g9698, g4725, g9964, g9954, g5523, g8550,
         g8402, g8845, g8611, g2081, g6359, g11586, g11007, g5147, g5104,
         g5099, g4821, g5919, g5499, g4389, g3529, g6416, g3497, g4990, g9619,
         g9010, I6630, g6047, g9652, g10505, g10469, g9843, g9711, g9519,
         g5273, g11465, g4348, g11237, g9834, g9731, g6654, g5444, g3714,
         g11285, g9598, g8097, g8726, g6880, g4816, g3287, g10759, g9938,
         g9917, g10758, g10652, g9909, g9891, g7127, g6663, g11165, g6328,
         g8401, g11006, g5125, g4865, g4715, g4604, g2325, g5513, g11222,
         g6554, g7732, g9586, g5178, g4401, g4104, g4584, g7472, g11253, g9860,
         g8703, g11600, g9645, g11236, g4162, g3106, g6090, g9691, g11316,
         g11175, g8068, g9607, g9962, g9952, g6348, g9659, g9358, I6316, I6317,
         g4486, g9587, g8995, g5632, g8965, g4881, g11209, g8848, g8715, g4070,
         g3263, g6463, g8699, g7820, g11021, g5917, g6619, g6318, g6872,
         g11201, g10514, g10489, g4006, g9853, g11274, g8119, g9420, g5233,
         g7092, g6549, g11464, g4487, g2939, g7060, g6739, g5725, g11615,
         g2544, g11252, g5532, g11153, g3771, g9905, g9872, g9680, g7739,
         g6321, g8386, g8975, g2306, g6625, g7937, g8303, g8170, g5706, g2756,
         g8821, g8643, g10946, g5225, g4169, g5029, g11164, g4007, g4059,
         g4868, g5675, g4718, g10682, g6687, g7704, g4261, g3422, g5745, g8387,
         g7954, g11283, g8461, g8298, g10760, g11480, g6626, g8756, g6341,
         g10506, g9648, g7453, g5995, g6645, g5707, g7548, g11091, g11174,
         g8403, g8841, g8605, g6879, g8763, g4502, g9839, g9702, g9742, g6358,
         g5841, g5575, g8107, g10240, g11192, g9618, g5539, g8416, g9693,
         g11553, g7557, g5268, g9107, g10633, g7894, g8654, g9621, g6794,
         g5819, g4883, g3412, g7661, g2800, g3389, g3268, g9908, g3429, g6628,
         g5470, g7526, g2204, g5025, g6204, g4921, g4048, g8935, g2525, g9593,
         g4827, g10701, g10777, g10733, g8130, g9965, g9955, g3684, g11213,
         g5006, g9933, g9912, g8554, g8407, g9641, g6323, g10766, g10646,
         g6666, g4994, g5103, g11592, g3717, g6875, g9658, g6530, g6207, g8199,
         g7265, g9835, g9735, g6655, g3875, g7970, g7384, g5491, g8949, g11152,
         g9611, g6410, g2804, g10451, g4397, g7224, g5398, g5602, g6884, g8698,
         g8964, g11413, g4950, g5535, g7277, g6772, g8463, g8301, g2511,
         g10728, g6618, g6235, g6355, g4723, g3626, g8720, g6693, g11020,
         g11583, g8118, g8167, g7892, g8652, g5721, g10367, g10362, g9901,
         g6792, g11282, g7945, g11302, g11105, g3634, g8598, g8471, g7140,
         g9600, g9864, g11613, g5188, g7435, g7876, g4058, g6776, g5809,
         g10301, g4505, g9623, g10739, g11027, g10738, g8687, g8558, g6360,
         g9871, g5108, g11248, g4992, g11552, g9651, g11204, g7824, g5115,
         g8710, g7102, g9384, g2561, g9838, g9700, g9754, g3718, g10661,
         g10594, g11321, g8879, g7621, g8962, g10715, g2272, g8659, g9643,
         g8957, g5538, g4000, g4126, g4400, g4088, I5886, I5887, g6238, g10727,
         g8174, g5067, g5418, g10297, g6353, g11026, g11212, g6744, g4828,
         g10671, g4383, g2517, g5256, g4297, g4220, g8380, g8252, g7071, g9613,
         g8933, g5181, g7948, g11149, g9862, g11387, g7955, g4161, g11148,
         g2321, g9712, g8931, g11097, g3819, g11104, g2963, g6092, g4999,
         g7409, g4976, g6858, g4103, I6309, g6580, g5944, g5631, g9414, g9660,
         g9946, g9926, I6331, g9903, g9885, g9673, g10625, g6623, g11228,
         g11011, g6889, g7523, g7822, g8123, g11582, g4316, g3400, g10969,
         g3625, g5041, g9335, g9831, g9727, g9422, g8648, g4588, g8511, g8875,
         g5168, g7895, g7503, g8655, g3396, g4914, g9947, g9927, g5772, g5531,
         g5036, g10503, g8010, g7738, g8410, g6231, g5608, g10581, g10450,
         g10364, g2132, g2379, g4820, g9653, g10818, g8172, g10429, g5074,
         g9869, g10741, g10635, g8693, g5480, g4581, g3766, g2981, g8555,
         g8409, g9364, g8994, g11299, g6592, g7958, g4995, g4079, g2264, g2160,
         g3257, I6310, g5000, g3301, I5084, g9412, g9389, g10706, g10567,
         g10366, g10447, g10446, g10533, g5220, g10624, g10300, g5023, g4432,
         g4053, g7596, g5588, g6074, g9963, g9953, g3772, g3089, g5051, g8724,
         g4157, g9707, g8878, g10763, g10639, g6777, g8109, g7898, g7511,
         g11271, g11461, g5732, g11145, g11031, g9865, g9715, g9604, g8799,
         g8647, g11198, g6873, g6632, g6095, g9833, g9729, g6102, g7819,
         g11280, g7088, g9584, g9896, g8209, g6752, g11161, g8947, g5681,
         g7951, g9419, g5533, g8936, g10670, g11087, g4949, g6364, g5851,
         g7825, g10667, g7136, g6532, g9385, g9897, g9425, g3383, g5601, g7943,
         g11171, I6631, g7230, g6064, g4952, g8736, g6787, g8968, g10306,
         g11459, g11458, g5739, g7496, g4986, g11010, g5187, g3999, g8175,
         g8722, g5590, g7891, g7471, g8651, g5479, g11599, g6684, g6745, g6639,
         g3696, g4503, g6791, g8180, g4224, g5501, g8838, g8602, g10666,
         g11158, g9602, g5704, g4617, g3879, g9868, g11295, g11144, g9718,
         g3434, g4987, g6098, g9582, g3533, g8104, g9415, g8499, g8377, g9664,
         g2534, g8754, g9413, g6162, g3584, g4991, g6362, g5846, g10685,
         g11023, g7598, g11224, g11571, g4959, g5626, g9940, g9920, g4876,
         g6730, g9689, g10762, g6070, g9428, g9430, g8927, g7068, g8014, g7740,
         g11278, g5782, g9910, g4236, g11559, g9609, g11558, g6087, g4877,
         g10751, g10772, g10655, g8135, g11544, g5084, g8382, g10230, g7241,
         g3942, g10638, g4064, g9365, g9861, g9738, g9579, g8749, g11255,
         g11189, g10510, g2917, g11188, g9846, g7818, g11460, g11030, g11093,
         g7893, g7478, g8653, g10442, g6535, g8102, I5085, g3912, g7186, g4489,
         g9662, g9418, g11218, g10746, g10643, g7125, g7821, g6246, g8963,
         g7533, g10237, g7939, g8786, g8638, g10684, g11455, g8364, g2990,
         g9847, g7584, g5617, g5981, g5789, g4009, g11277, g6940, g6472, g7061,
         g6760, g11595, g5771, g8553, g8405, g4836, g5547, g4967, g6671, g7200,
         g7046, g4229, g8389, g6430, g8706, g4993, g6247, g11170, g7145, g5738,
         g3998, g6741, g11167, g11194, g11589, g4431, g7536, g9585, g2957,
         g11588, g5690, g6883, g4837, g8791, g8641, g6217, g11022, g5915,
         g4168, g8759, g5110, g11254, g7567, g4392, g3273, g9856, g9411, g5002,
         g11101, g11177, g11560, g8098, g3970, g4941, g6662, g7935, g6067,
         g9863, g9740, g6994, g6758, g4252, g11166, g7130, g11009, g5179,
         g7542, g11008, g5171, g3516, g7573, g3987, g11555, g9857, g9734,
         g9569, g8728, g8730, g8185, g8385, g7902, g4073, g8070, g5731, g11238,
         g8470, g8308, g5489, g3991, g7823, g4069, g11176, g11092, g11154,
         g9608, g11637, g2091, g8406, g5254, g8612, g9588, g8801, g8742, g7063,
         g10303, g5009, g9665, g8748, g11215, g10750, g5769, g3818, g8755,
         g6673, g7720, g4609, g7547, g7971, g11288, g7599, g6058, g6743, g4106,
         g6890, g7549, g7269, g8169, g11304, g9944, g9924, g7592, g8718, g8616,
         g9316, g7625, g8793, g8644, g2940, g11624, g10949, g2947, g4870,
         g3563, g10948, g2223, g8246, g7846, g5788, g4008, g9596, g5249,
         g11585, g4972, g11554, g7096, g10673, g4806, g2493, g9936, g9915,
         g2910, g9317, g10933, g10853, g8388, g8177, g7141, g10508, g4230,
         g10634, g9601, g9192, g6326, g7710, g8028, g7375, g5640, g5031, g4550,
         g7879, g7962, g9597, g5005, g6423, g8108, g5911, g3322, g9937, g9916,
         g9840, g9704, g9747, g10723, g8217, g11013, g5209, g9390, g11214,
         g6327, g5796, g5473, g6346, g5038, g6633, g11005, g5119, g8365, g7558,
         g4481, g4097, g7588, g4497, g9942, g9922, g6696, g10731, g5118,
         g10665, g8827, g8552, g5540, g4960, g8846, g8615, g5983, g6240, g7931,
         g11100, g11235, g5199, g6316, g7515, g5781, g8018, g7742, g2950,
         g5510, g6347, g9357, g11407, g10743, g5259, g5694, g10769, g11584,
         g4932, g10768, g10649, g4068, g6317, g5215, g4276, g4866, g6775,
         g10662, g8101, g5825, g3204, g5318, g7884, g7457, g3974, g9949, g9929,
         g10778, g7524, g6079, g7235, g9603, g9850, g9726, g9560, g7988, g5228,
         g5587, g5934, g8168, g9583, g10672, g8627, g8309, g10449, g10420,
         g11273, g8734, g5913, g4572, g6363, g11463, g8074, g8474, g8383,
         g11234, g4483, g11491, g5097, g5726, g5497, g7933, g9617, g9906,
         g9873, g9683, g11012, g5196, g7050, g10971, g10849, g8400, g4345,
         g9945, g9925, g7271, g5028, g9709, g4223, g10716, g10497, g11247,
         g6661, g11173, g6075, g8023, g7367, g9907, g9888, g9686, g10582,
         g5746, g9959, g9950, g7674, g9690, g5703, g4522, g4115, g7075, g10627,
         g4047, g2944, g6646, g7132, g11029, g7572, g8127, g7209, g11028,
         g10742, g8880, g10681, g9663, g5349, g8732, g3807, g8753, g5848,
         g3860, g8508, g8411, g8072, g5699, g11240, g6616, g6105, g10690,
         g7582, g9590, g4128, g6404, g6647, g10504, g9657, g4542, g5524, g9899,
         g7736, g10626, g6320, g7623, g10299, g7889, g10298, g8413, g3979,
         g5211, g4512, g7722, g9844, g9714, g9522, g4823, g5993, g5026, g8705,
         g10737, g10232, g6771, g5170, g8117, g9966, g9956, g5280, g7139,
         g11099, g6892, g9705, g10512, g11098, g8628, g5544, g11272, g5483,
         g9948, g9928, g4063, g11462, g6738, g7593, g11032, g10445, g8882,
         g10316, g5756, g4720, g9409, g8929, g6876, g4989, g9836, g9737, g6061,
         g8268, g6465, g5003, g9967, g9957, g5145, g4834, g4971, g10753, g5695,
         g7613, g10736, g11220, g7444, g4670, g4253, g8163, g7960, g10764,
         g5757, g10365, g8032, g7385, g11591, g2988, g7583, g11147, g5522,
         g9837, g9697, g9751, g9620, g11151, g11172, g7885, g5595, g5537,
         g9842, g9708, g9516, g4141, g4341, g7679, g7378, g5612, g3939, g7135,
         g10970, g11025, g9854, g9730, g9566, g7182, g9941, g9921, g6194,
         g4962, g4358, g8683, g4803, g8549, g5224, g8778, g11281, g8735,
         g11146, g3904, g2948, g8075, g9829, g9723, g7184, g11246, g6350,
         g5837, g5902, g2555, g6438, g5512, g5090, g7719, g3695, g7587, g9610,
         g3536, g8881, g4559, g10561, g10549, g5698, g11226, g10295, g5260,
         g10680, g11551, g11538, g9849, g5279, g8404, g5720, g8764, g11318,
         g11297, g9898, g9510, g7963, g9759, g9803, g6124, I14585, I5600,
         g9489, g3107, g2167, g9362, I14866, g4997, g10291, g9669, g6122,
         g9509, g5227, I15054, g5555, g10376, g8249, I15210, g9882, I5805,
         g2102, g2099, g2096, g2088, I15039, g8259, g10805, I15214, I15215,
         g8322, g9750, g8248, g8154, I6351, g2405, g2389, g2380, g2372, I16427,
         I14776, g4052, g2862, g2515, I14858, I15209, g2528, g2522, g9515,
         g3118, g2180, I5571, g2514, I5599, g9528, I5629, g2315, I5363, g8159,
         g10521, I16148, I16149, g8417, I14855, I15205, g9878, I15051, g9615,
         g8823, g8148, g2863, g2516, g9511, g9654, I15224, I15225, g8253,
         g9416, I15171, I15172, g9410, I15204, I14596, g9655, g10472, g10470,
         g10468, g10467, g10386, g10384, g10476, g10474, g8158, g9656, g9746,
         I5357, g9758, I5626, I15057, I15219, I15220, g9616, I14862, g2521,
         I14751, g9591, g9757, g9815, I14835, I16161, g10479, g10478, g10477,
         g10475, g2353, g9776, I5804, I15199, g8153, g9881, g9426, g9423,
         g8262, g2499, I5570, I14607, g9388, g10807, I16160, g10394, g10392,
         g10482, g10481, I15042, g9589, g9667, I14827, g9779, g9391, g2309,
         I5358, I15177, g9876, g9421, g5186, I6350, g8162, I14779, g2305,
         I5351, I5352, I15176, g9879, g10562, g9606, I14822, I15200, g9880,
         I14582, g8247, I5576, g4476, g2538, I5649, g9605, g9781, g9363,
         I14831, g8263, g9361, g5780, I15048, g9647, g9817, I14602, I15033,
         g2445, g2437, g2433, g2419, I5366, g9506, g8161, g2316, g4675, g9387,
         I15045, g9808, g2501, g9877, g10529, g9874, g8157, g6899, g9646,
         g2111, g2109, g2106, g2104, I5612, I5613, I5593, I5591, g8970, g8839,
         I10519, I11279, I11278, g3978, I5264, I5263, I8640, g4278, I6761,
         g2943, I6760, I17400, g11418, g11416, I5450, I5449, I16060, g10372,
         I16058, I6746, g2938, I11975, I11973, I12136, I11937, I11935, g2959,
         I6167, I6168, I5878, g2120, g2115, I5619, I5620, g5552, I6468, I6467,
         I8796, g4672, I8795, I15891, I15892, I5611, g8738, I6716, I6714,
         I7685, g3460, I7683, I12108, I12106, I6747, g2236, I5230, I5231,
         I12075, I12076, I15870, g10358, I16067, I16065, I7562, I13531, I13529,
         I8797, I17584, I11936, I15257, I15256, I13505, I13506, g8824, g8502,
         g8501, I6186, g11496, I17504, I17505, I16001, I15999, I6125, g2215,
         I6124, I11909, I11907, I12040, I12038, I13909, I13907, I6771, I6772,
         I11908, I16008, I16009, I13908, I7034, I7035, I8650, I9947, I9948,
         I16066, g10428, I6144, I6145, I11242, I11241, I15993, I15994, I6187,
         g6027, I5500, I11974, I12062, I12060, I8771, I8772, I5184, I13293,
         I6200, I6199, I13265, I5024, I5023, I7863, I13991, I13992, I13660,
         I13661, I6143, I13990, I11510, I11508, g5034, I5229, I12047, I12045,
         I10771, I10769, I16045, I16046, I12061, I5104, I13530, I6447, I4956,
         I4954, I8481, g3530, I8479, I8739, I8740, I6880, I6879, I15431,
         I15430, I12020, I12019, I16331, I16332, I16469, I16467, I5014, I5013,
         I13523, I13521, I16039, I16037, I16468, I12046, I16038, g10427, I8676,
         g4374, I12113, I8761, g4616, g10422, I15992, I5036, I5034, I14263,
         g8843, I13249, I13250, I5135, I5485, I5486, I7033, I15443, I15441,
         I6166, I8624, g4267, I16015, g10425, I8677, I8576, g4234, I8575,
         I14613, g9204, I14612, I8716, g4601, I8715, I6715, I13514, I13515,
         I12003, I12002, g2177, I5127, I5128, I8577, I17395, g11414, I17393,
         I11280, I5265, I6989, I6988, I13274, I13272, I10507, I5164, I14443,
         I14444, I9559, I9557, I5592, I13077, I13078, I8717, I5296, I5295,
         I8625, I8626, I4911, I4912, I16000, g10423, I5371, I5185, I5186,
         I5675, I8544, g4218, I8543, I10520, I10521, I5297, I13537, I13283,
         g4749, I11982, I11980, I8514, g4873, I8513, I13091, I13089, I6126,
         I15908, g10302, I15906, I8763, g8825, g8506, I16007, g10424, I5865,
         g2107, g2105, I5604, I5517, I5518, I6111, I6109, I4929, I4930, I13522,
         I10770, I5539, I5538, I17394, g11415, I13553, I13552, I8642, I17296,
         I17297, I14278, I14279, I4910, I6794, I6792, I5484, I15442, I10931,
         I10932, I8779, I8780, g2354, I15615, g10043, g10153, I17281, I5470,
         I5468, I11509, I5025, I14272, I14270, I6208, I6209, I17290, I17288,
         I7563, I7564, I5006, I5005, I12128, I12126, I5105, I6323, I6322,
         I12093, I12094, I6666, g2776, I6664, g3623, I6762, I5373, I8529,
         I8527, I5283, I5282, I7224, I7223, I5007, I5459, I17295, I5015,
         I14264, I14265, I16073, I16072, g3205, I8652, I9558, I5203, I5202,
         I6806, I6807, I6469, I12145, I12143, I12127, I13302, I13300, I5502,
         I9574, I6448, I6449, I8670, I8669, I15453, I15451, I7876, I7875,
         I14203, I14202, I15607, g10149, g10144, I5324, I5325, I8738, g10434,
         g5859, I8606, I8604, I12087, I12085, I13248, I4979, I4980, I12069,
         I12067, g8942, I12068, I17503, I7877, I5165, I6289, I6287, I6777,
         I8562, I8563, I15890, I13090, g8006, g11474, I17460, I17461, I13513,
         I4986, I4987, I5204, I13504, I6207, I12086, I8545, I8180, I8178,
         I8591, I8589, I10930, I17402, I13294, I13295, I12144, g8757, g2961,
         I14211, I14209, I8515, I5316, I5317, I9946, I8750, g4613, I5605,
         I14204, I16051, g10371, g10373, g10360, g6037, I13858, I13859, I15872,
         I8528, g4879, I13901, I13902, g8542, I6838, I6836, I17307, I17305,
         g4538, I15452, I13857, I13765, I8671, g10370, I16044, g10363, g5360,
         I5106, I8804, g4677, I8803, I16016, I16017, I17487, I17485, I4995,
         I12092, I8678, I5126, I5372, I17306, I11995, I7225, I11261, g8545,
         I6110, I4942, I4941, I15899, I15900, g5527, g10443, g5350, I16081,
         g10374, I16079, I8641, I6178, I6176, I12074, I5451, I7322, I7323,
         I6288, I8179, I6805, I17486, I4928, g10286, I16330, I9575, I13887,
         I13886, I8787, I8788, I5315, g10285, I13869, I13867, I13868, I13259,
         I13258, g3261, I16074, I5136, I5137, I5460, I5461, I8605, I6770,
         g11449, I17401, g11448, I15717, g10231, I15716, I14210, I17569,
         I17567, I13878, I13876, I5606, I14442, I11996, I11997, I14277, I17568,
         I7321, I6990, g8847, I9006, I4985, I8651, I13545, I13544, I13894,
         I13895, I6138, I6136, I13076, g2205, I13260, I5501, I17586, I13900,
         I6201, I14217, g8826, I14216, I9007, I13561, I13559, g10229, I17493,
         I17492, I12215, I12214, I11262, I11263, I6225, I6226, I13309, I13307,
         I5676, I5677, I6826, I6827, I13308, g8190, g2792, I5879, I5880, g3061,
         I17585, I6881, I12138, I8729, g4605, I8728, I15871, I5866, I5867,
         I6793, I6487, I16080, I13893, I12115, I6748, I6224, I8805, I15880,
         I15878, I16031, I16030, I14271, I13267, I15616, I15617, I4966, I4964,
         I8752, I15432, g10438, g6032, g3011, I8480, I16087, I16086, g3734,
         I14218, I4955, I8786, g4639, g10480, I11915, I11914, I8770, g4619,
         I5516, g8541, I6188, I5892, I5891, I13766, I13767, I15258, I13266,
         I6825, I17283, g5277, I5035, g10375, I15879, g10359, I12114, I12107,
         g2500, g10430, g5999, I13285, I13877, g2795, I5893, I13560, g4259,
         I5166, I14614, I4965, I4943, I16023, g10426, I16059, g8737, I9576,
         I16052, I16053, I12004, g5573, I6837, I8730, I4978, I6177, I17051,
         I7864, I7865, I6665, I12216, I13554, g10368, I13284, I6137, I5529,
         I5530, I17282, I5618, I8664, I8662, I11916, g7717, I4972, I4971,
         I13273, I10509, I10508, I6778, I6779, I5469, g4251, I13546, I4996,
         I4997, I13539, I16032, I5323, I13538, I5540, I8778, g4286, I17052,
         I17053, g10287, I15898, g7978, g4227, I8561, I8762, I8751, I15907,
         I4973, I16024, I16025, g4455, I5342, I5341, I12137, g10483, I16088,
         I17289, g4630, I15609, I15608, g10436, g6023, I17459, I13301, I11981,
         I8663, I15718, I5284, g4607, g8840, g10441, g5345, g10432, g5938,
         I12021, I6489, I5528, I13659, I5343, I12039, I9008, I6488, I13888,
         I17494, I7684, g3221, I6324, I8590, I11243, g10324, g10239, g4974,
         g10322, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, g5816, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1301, n1302, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1388, n1389, n1390, n1391, n1392;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4207 = g1200;
  assign g4208 = g1203;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g8061 = g872;
  assign g5101 = g872;
  assign g8062 = g873;
  assign g5105 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g4177 = g774;
  assign g4180 = g786;
  assign g3007 = g878;
  assign g2602 = g587;
  assign g2609 = g583;
  assign g4173 = g758;
  assign g2986 = g883;
  assign g2605 = g579;
  assign g4175 = g766;
  assign g2603 = g588;
  assign g2606 = g580;
  assign g2612 = g586;
  assign g3069 = g1206;
  assign g4178 = g778;
  assign g4176 = g770;
  assign g2648 = g865;
  assign g4179 = g782;
  assign g2601 = g578;
  assign g4174 = g762;
  assign g2604 = g589;
  assign g4172 = g754;
  assign g4181 = g790;
  assign g2608 = g582;
  assign g2610 = g584;
  assign g2607 = g581;
  assign g2611 = g585;
  assign g8565 = g3435;
  assign g6949 = g3435;
  assign g10459 = g10408;
  assign g10377 = g10336;
  assign g8561 = g3399;
  assign g6920 = g3399;
  assign g8331 = g8226;
  assign g8982 = g8814;
  assign g10465 = g10417;
  assign g9961 = g9931;
  assign g8349 = g8241;
  assign g10457 = g10405;
  assign g8323 = g8214;
  assign g8352 = g8187;
  assign g8564 = g3431;
  assign g6942 = g3431;
  assign g10801 = g10712;
  assign g4171 = g2791;
  assign g10461 = g10411;
  assign g8313 = g8203;
  assign g10463 = g10414;
  assign g5659 = g3418;
  assign g8984 = g8816;
  assign g9451 = g9088;
  assign g10628 = g10515;
  assign g8983 = g8815;
  assign g11206 = g10583;
  assign g8563 = g3425;
  assign g6932 = g3425;
  assign g11163 = g10779;
  assign g8566 = g3438;
  assign g6955 = g3438;
  assign g8562 = g3414;
  assign g6926 = g3414;
  assign g8980 = g8812;
  assign g10455 = g10402;
  assign g8328 = g8221;
  assign g8347 = g8200;
  assign g8979 = g8811;
  assign g11489 = g11425;
  assign g8985 = g8818;
  assign g8340 = g8236;
  assign g10379 = g10339;
  assign g8316 = g8206;
  assign g8976 = g8817;
  assign g8978 = g8810;
  assign g8335 = g8230;
  assign g6842 = g5287;
  assign g8986 = g8819;
  assign g5658 = g3407;
  assign g8977 = g8806;
  assign g8981 = g8813;
  assign g8318 = g8210;
  assign g8271 = g5816;

  dff_0 DFF_0 ( .clk(CK), .q(g1289), .d(g4556) );
  dff_533 DFF_1 ( .clk(CK), .q(g1882), .d(g8943) );
  dff_532 DFF_2 ( .clk(CK), .q(g312), .d(g255) );
  dff_531 DFF_3 ( .clk(CK), .q(g452), .d(g11257) );
  dff_530 DFF_4 ( .clk(CK), .q(g123), .d(g7032) );
  dff_529 DFF_5 ( .clk(CK), .q(g207), .d(g6830) );
  dff_528 DFF_6 ( .clk(CK), .q(g713), .d(g8920) );
  dff_527 DFF_7 ( .clk(CK), .q(g1153), .d(g4340) );
  dff_526 DFF_8 ( .clk(CK), .q(g1209), .d(g10732) );
  dff_525 DFF_9 ( .clk(CK), .q(g1744), .d(g4239) );
  dff_524 DFF_10 ( .clk(CK), .q(g1558), .d(g6538) );
  dff_523 DFF_11 ( .clk(CK), .q(g695), .d(g8887) );
  dff_522 DFF_12 ( .clk(CK), .q(g461), .d(g11372) );
  dff_521 DFF_13 ( .clk(CK), .q(g940), .d(g8260) );
  dff_520 DFF_14 ( .clk(CK), .q(g976), .d(g11391) );
  dff_519 DFF_15 ( .clk(CK), .q(g709), .d(g8432) );
  dff_518 DFF_16 ( .clk(CK), .q(g1092), .d(g6088) );
  dff_517 DFF_17 ( .clk(CK), .q(g1574), .d(g6478) );
  dff_516 DFF_18 ( .clk(CK), .q(g1864), .d(g6795) );
  dff_515 DFF_19 ( .clk(CK), .q(g369), .d(g11320) );
  dff_514 DFF_20 ( .clk(CK), .q(g1580), .d(g6500) );
  dff_513 DFF_21 ( .clk(CK), .q(g1736), .d(g5392) );
  dff_512 DFF_22 ( .clk(CK), .q(g39), .d(g10663) );
  dff_511 DFF_23 ( .clk(CK), .q(g1651), .d(g10782) );
  dff_510 DFF_24 ( .clk(CK), .q(g1424), .d(g6216) );
  dff_509 DFF_25 ( .clk(CK), .q(g1737), .d(g1736) );
  dff_508 DFF_26 ( .clk(CK), .q(g1672), .d(g10858) );
  dff_507 DFF_27 ( .clk(CK), .q(g1077), .d(g5914) );
  dff_506 DFF_28 ( .clk(CK), .q(g1231), .d(g7590) );
  dff_505 DFF_29 ( .clk(CK), .q(g4), .d(g6656) );
  dff_504 DFF_30 ( .clk(CK), .q(g774), .d(g6728) );
  dff_503 DFF_31 ( .clk(CK), .q(g1104), .d(g5126) );
  dff_502 DFF_32 ( .clk(CK), .q(g1304), .d(g7290) );
  dff_501 DFF_33 ( .clk(CK), .q(g243), .d(g6841) );
  dff_500 DFF_34 ( .clk(CK), .q(g1499), .d(g8041) );
  dff_499 DFF_35 ( .clk(CK), .q(g1044), .d(g7106) );
  dff_498 DFF_36 ( .clk(CK), .q(g1444), .d(g8766) );
  dff_497 DFF_37 ( .clk(CK), .q(g757), .d(g10788) );
  dff_496 DFF_38 ( .clk(CK), .q(g786), .d(g8019) );
  dff_495 DFF_39 ( .clk(CK), .q(g1543), .d(g6545) );
  dff_494 DFF_40 ( .clk(CK), .q(g552), .d(g10856) );
  dff_493 DFF_41 ( .clk(CK), .q(g315), .d(g256) );
  dff_492 DFF_42 ( .clk(CK), .q(g1534), .d(g6533) );
  dff_491 DFF_43 ( .clk(CK), .q(g622), .d(g8820) );
  dff_490 DFF_44 ( .clk(CK), .q(g1927), .d(g8941) );
  dff_489 DFF_45 ( .clk(CK), .q(g1660), .d(g10859) );
  dff_488 DFF_46 ( .clk(CK), .q(g278), .d(g6922) );
  dff_487 DFF_47 ( .clk(CK), .q(g1436), .d(g8772) );
  dff_486 DFF_48 ( .clk(CK), .q(g718), .d(g8433) );
  dff_485 DFF_49 ( .clk(CK), .q(g76), .d(g6526) );
  dff_484 DFF_50 ( .clk(CK), .q(g554), .d(g10793) );
  dff_483 DFF_51 ( .clk(CK), .q(g496), .d(g11333) );
  dff_482 DFF_52 ( .clk(CK), .q(g981), .d(g11392) );
  dff_481 DFF_53 ( .clk(CK), .q(g878), .d(g3506) );
  dff_480 DFF_54 ( .clk(CK), .q(g590), .d(g1713) );
  dff_479 DFF_55 ( .clk(CK), .q(g829), .d(g794) );
  dff_478 DFF_56 ( .clk(CK), .q(g1095), .d(g6093) );
  dff_477 DFF_57 ( .clk(CK), .q(g704), .d(g8889) );
  dff_476 DFF_58 ( .clk(CK), .q(g1265), .d(g7302) );
  dff_475 DFF_59 ( .clk(CK), .q(g1786), .d(g6525) );
  dff_474 DFF_60 ( .clk(CK), .q(g682), .d(g8429) );
  dff_473 DFF_61 ( .clk(CK), .q(g1296), .d(g7292) );
  dff_472 DFF_62 ( .clk(CK), .q(g587), .d(g104) );
  dff_471 DFF_63 ( .clk(CK), .q(g52), .d(g6621) );
  dff_470 DFF_64 ( .clk(CK), .q(g646), .d(g7134) );
  dff_469 DFF_65 ( .clk(CK), .q(g327), .d(g260) );
  dff_468 DFF_66 ( .clk(CK), .q(g1389), .d(g6333) );
  dff_467 DFF_67 ( .clk(CK), .q(g1371), .d(g6826) );
  dff_466 DFF_68 ( .clk(CK), .q(g1956), .d(g1955) );
  dff_465 DFF_69 ( .clk(CK), .q(g1675), .d(g10860) );
  dff_464 DFF_70 ( .clk(CK), .q(g354), .d(g11483) );
  dff_463 DFF_71 ( .clk(CK), .q(g113), .d(g6392) );
  dff_462 DFF_72 ( .clk(CK), .q(g639), .d(g7626) );
  dff_461 DFF_73 ( .clk(CK), .q(g1684), .d(g10866) );
  dff_460 DFF_74 ( .clk(CK), .q(g1639), .d(g8193) );
  dff_459 DFF_75 ( .clk(CK), .q(g1791), .d(g6983) );
  dff_458 DFF_76 ( .clk(CK), .q(g248), .d(g6839) );
  dff_457 DFF_77 ( .clk(CK), .q(g1707), .d(g4076) );
  dff_456 DFF_78 ( .clk(CK), .q(g1759), .d(g4293) );
  dff_455 DFF_79 ( .clk(CK), .q(g351), .d(g11482) );
  dff_454 DFF_80 ( .clk(CK), .q(g1957), .d(g1956) );
  dff_453 DFF_81 ( .clk(CK), .q(g1604), .d(g6507) );
  dff_452 DFF_82 ( .clk(CK), .q(g1098), .d(g6096) );
  dff_451 DFF_83 ( .clk(CK), .q(g932), .d(g8250) );
  dff_450 DFF_84 ( .clk(CK), .q(g126), .d(g2807) );
  dff_449 DFF_85 ( .clk(CK), .q(g1896), .d(g8282) );
  dff_448 DFF_86 ( .clk(CK), .q(g736), .d(g8435) );
  dff_447 DFF_87 ( .clk(CK), .q(g1019), .d(g6924) );
  dff_446 DFF_88 ( .clk(CK), .q(g1362), .d(g6819) );
  dff_445 DFF_89 ( .clk(CK), .q(g745), .d(g746) );
  dff_444 DFF_90 ( .clk(CK), .q(g1419), .d(g6244) );
  dff_443 DFF_91 ( .clk(CK), .q(g58), .d(g6627) );
  dff_442 DFF_92 ( .clk(CK), .q(g32), .d(g11286) );
  dff_441 DFF_93 ( .clk(CK), .q(g876), .d(g878) );
  dff_440 DFF_94 ( .clk(CK), .q(g1086), .d(g6071) );
  dff_439 DFF_95 ( .clk(CK), .q(g1486), .d(g8046) );
  dff_438 DFF_96 ( .clk(CK), .q(g1730), .d(g10707) );
  dff_437 DFF_97 ( .clk(CK), .q(g1504), .d(g6198) );
  dff_436 DFF_98 ( .clk(CK), .q(g1470), .d(g8051) );
  dff_435 DFF_99 ( .clk(CK), .q(g822), .d(g8024) );
  dff_434 DFF_100 ( .clk(CK), .q(g583), .d(g29) );
  dff_433 DFF_101 ( .clk(CK), .q(g1678), .d(g10862) );
  dff_432 DFF_102 ( .clk(CK), .q(g174), .d(g8050) );
  dff_431 DFF_103 ( .clk(CK), .q(g1766), .d(g7133) );
  dff_430 DFF_104 ( .clk(CK), .q(g1801), .d(g7930) );
  dff_429 DFF_105 ( .clk(CK), .q(g186), .d(g6832) );
  dff_428 DFF_106 ( .clk(CK), .q(g959), .d(g11308) );
  dff_427 DFF_107 ( .clk(CK), .q(g1169), .d(g5189) );
  dff_426 DFF_108 ( .clk(CK), .q(g1007), .d(g6918) );
  dff_425 DFF_109 ( .clk(CK), .q(g1407), .d(g8769) );
  dff_424 DFF_110 ( .clk(CK), .q(g1059), .d(g7236) );
  dff_423 DFF_111 ( .clk(CK), .q(g1868), .d(g6909) );
  dff_422 DFF_112 ( .clk(CK), .q(g758), .d(g4940) );
  dff_421 DFF_113 ( .clk(CK), .q(g1718), .d(g5404) );
  dff_420 DFF_114 ( .clk(CK), .q(g396), .d(g11265) );
  dff_419 DFF_115 ( .clk(CK), .q(g1015), .d(g6930) );
  dff_418 DFF_116 ( .clk(CK), .q(g38), .d(g10726) );
  dff_417 DFF_117 ( .clk(CK), .q(g632), .d(g4891) );
  dff_416 DFF_118 ( .clk(CK), .q(g1415), .d(g6224) );
  dff_415 DFF_119 ( .clk(CK), .q(g1227), .d(g7586) );
  dff_414 DFF_120 ( .clk(CK), .q(g1721), .d(g10770) );
  dff_413 DFF_121 ( .clk(CK), .q(g882), .d(g883) );
  dff_412 DFF_122 ( .clk(CK), .q(g16), .d(g3524) );
  dff_411 DFF_123 ( .clk(CK), .q(g284), .d(g6934) );
  dff_410 DFF_124 ( .clk(CK), .q(g426), .d(g11256) );
  dff_409 DFF_125 ( .clk(CK), .q(g219), .d(g6824) );
  dff_408 DFF_126 ( .clk(CK), .q(g1216), .d(g1360) );
  dff_407 DFF_127 ( .clk(CK), .q(g806), .d(g6126) );
  dff_406 DFF_128 ( .clk(CK), .q(g1428), .d(g8767) );
  dff_405 DFF_129 ( .clk(CK), .q(g579), .d(g102) );
  dff_404 DFF_130 ( .clk(CK), .q(g1564), .d(g6546) );
  dff_403 DFF_131 ( .clk(CK), .q(g1741), .d(g4238) );
  dff_402 DFF_132 ( .clk(CK), .q(g225), .d(g6823) );
  dff_401 DFF_133 ( .clk(CK), .q(g281), .d(g6928) );
  dff_400 DFF_134 ( .clk(CK), .q(g1308), .d(g11602) );
  dff_399 DFF_135 ( .clk(CK), .q(g611), .d(g9721) );
  dff_398 DFF_136 ( .clk(CK), .q(g631), .d(g4890) );
  dff_397 DFF_137 ( .clk(CK), .q(g1217), .d(n1197) );
  dff_396 DFF_138 ( .clk(CK), .q(g1589), .d(g6524) );
  dff_395 DFF_139 ( .clk(CK), .q(g1466), .d(g8045) );
  dff_394 DFF_140 ( .clk(CK), .q(g1571), .d(g6469) );
  dff_393 DFF_141 ( .clk(CK), .q(g1861), .d(g6471) );
  dff_392 DFF_142 ( .clk(CK), .q(g1365), .d(g6821) );
  dff_391 DFF_143 ( .clk(CK), .q(g1448), .d(g11514) );
  dff_390 DFF_144 ( .clk(CK), .q(g1711), .d(g5403) );
  dff_389 DFF_145 ( .clk(CK), .q(g1133), .d(g4480) );
  dff_388 DFF_146 ( .clk(CK), .q(g1333), .d(g11610) );
  dff_387 DFF_147 ( .clk(CK), .q(g153), .d(g7843) );
  dff_386 DFF_148 ( .clk(CK), .q(g962), .d(g11310) );
  dff_385 DFF_149 ( .clk(CK), .q(g766), .d(g5536) );
  dff_384 DFF_150 ( .clk(CK), .q(g588), .d(g28) );
  dff_383 DFF_151 ( .clk(CK), .q(g486), .d(g11331) );
  dff_382 DFF_152 ( .clk(CK), .q(g471), .d(g11380) );
  dff_381 DFF_153 ( .clk(CK), .q(g1397), .d(g6838) );
  dff_380 DFF_154 ( .clk(CK), .q(g580), .d(g103) );
  dff_379 DFF_155 ( .clk(CK), .q(g1950), .d(g8288) );
  dff_378 DFF_156 ( .clk(CK), .q(g756), .d(g755) );
  dff_377 DFF_157 ( .clk(CK), .q(g635), .d(g4892) );
  dff_376 DFF_158 ( .clk(CK), .q(g1101), .d(g5390) );
  dff_375 DFF_159 ( .clk(CK), .q(g549), .d(g10855) );
  dff_374 DFF_160 ( .clk(CK), .q(g1041), .d(g7258) );
  dff_373 DFF_161 ( .clk(CK), .q(g105), .d(g10898) );
  dff_372 DFF_162 ( .clk(CK), .q(g1669), .d(g10865) );
  dff_371 DFF_163 ( .clk(CK), .q(g1368), .d(g6822) );
  dff_370 DFF_164 ( .clk(CK), .q(g1531), .d(g6528) );
  dff_369 DFF_165 ( .clk(CK), .q(g1458), .d(g6180) );
  dff_368 DFF_166 ( .clk(CK), .q(g572), .d(g10718) );
  dff_367 DFF_167 ( .clk(CK), .q(g1011), .d(g6912) );
  dff_366 DFF_168 ( .clk(CK), .q(g33), .d(g10719) );
  dff_365 DFF_169 ( .clk(CK), .q(g1411), .d(g6234) );
  dff_364 DFF_170 ( .clk(CK), .q(g1074), .d(g6099) );
  dff_363 DFF_171 ( .clk(CK), .q(g444), .d(g11259) );
  dff_362 DFF_172 ( .clk(CK), .q(g1474), .d(g8039) );
  dff_361 DFF_173 ( .clk(CK), .q(g1080), .d(g6059) );
  dff_360 DFF_174 ( .clk(CK), .q(g1713), .d(g5396) );
  dff_359 DFF_175 ( .clk(CK), .q(g333), .d(g262) );
  dff_358 DFF_176 ( .clk(CK), .q(g269), .d(g6906) );
  dff_357 DFF_177 ( .clk(CK), .q(g401), .d(g11266) );
  dff_356 DFF_178 ( .clk(CK), .q(g1857), .d(g11294) );
  dff_355 DFF_179 ( .clk(CK), .q(g9), .d(g5421) );
  dff_354 DFF_180 ( .clk(CK), .q(g664), .d(g8649) );
  dff_353 DFF_181 ( .clk(CK), .q(g965), .d(g11312) );
  dff_352 DFF_182 ( .clk(CK), .q(g1400), .d(g6840) );
  dff_351 DFF_183 ( .clk(CK), .q(g309), .d(g254) );
  dff_350 DFF_184 ( .clk(CK), .q(g814), .d(g7202) );
  dff_349 DFF_185 ( .clk(CK), .q(g231), .d(g6834) );
  dff_348 DFF_186 ( .clk(CK), .q(g557), .d(g10795) );
  dff_347 DFF_187 ( .clk(CK), .q(g586), .d(g103) );
  dff_346 DFF_188 ( .clk(CK), .q(g869), .d(g875) );
  dff_345 DFF_189 ( .clk(CK), .q(g1383), .d(g6831) );
  dff_344 DFF_190 ( .clk(CK), .q(g158), .d(g8060) );
  dff_343 DFF_191 ( .clk(CK), .q(g627), .d(g4893) );
  dff_342 DFF_192 ( .clk(CK), .q(g1023), .d(g7244) );
  dff_341 DFF_193 ( .clk(CK), .q(g259), .d(g6026) );
  dff_340 DFF_194 ( .clk(CK), .q(g1361), .d(g1206) );
  dff_339 DFF_195 ( .clk(CK), .q(g1327), .d(g11608) );
  dff_338 DFF_196 ( .clk(CK), .q(g654), .d(g7660) );
  dff_337 DFF_197 ( .clk(CK), .q(g293), .d(g6911) );
  dff_336 DFF_198 ( .clk(CK), .q(g1346), .d(g11640) );
  dff_335 DFF_199 ( .clk(CK), .q(g1633), .d(g8777) );
  dff_334 DFF_200 ( .clk(CK), .q(g1753), .d(g4274) );
  dff_333 DFF_201 ( .clk(CK), .q(g1508), .d(g6215) );
  dff_332 DFF_202 ( .clk(CK), .q(g1240), .d(g7297) );
  dff_331 DFF_203 ( .clk(CK), .q(g538), .d(g11326) );
  dff_330 DFF_204 ( .clk(CK), .q(g416), .d(g11269) );
  dff_329 DFF_205 ( .clk(CK), .q(g542), .d(g11325) );
  dff_328 DFF_206 ( .clk(CK), .q(g1681), .d(g10864) );
  dff_327 DFF_207 ( .clk(CK), .q(g374), .d(g11290) );
  dff_326 DFF_208 ( .clk(CK), .q(g563), .d(g10798) );
  dff_325 DFF_209 ( .clk(CK), .q(g1914), .d(g8284) );
  dff_324 DFF_210 ( .clk(CK), .q(g530), .d(g11328) );
  dff_323 DFF_211 ( .clk(CK), .q(g575), .d(g10800) );
  dff_322 DFF_212 ( .clk(CK), .q(g1936), .d(g8944) );
  dff_321 DFF_213 ( .clk(CK), .q(g55), .d(g7183) );
  dff_320 DFF_214 ( .clk(CK), .q(g1117), .d(g4465) );
  dff_319 DFF_215 ( .clk(CK), .q(g1317), .d(g1356) );
  dff_318 DFF_216 ( .clk(CK), .q(g357), .d(g11484) );
  dff_317 DFF_217 ( .clk(CK), .q(g386), .d(g11263) );
  dff_316 DFF_218 ( .clk(CK), .q(g1601), .d(g6501) );
  dff_315 DFF_219 ( .clk(CK), .q(g553), .d(g10857) );
  dff_314 DFF_220 ( .clk(CK), .q(g166), .d(g6757) );
  dff_313 DFF_221 ( .clk(CK), .q(g501), .d(g11334) );
  dff_312 DFF_222 ( .clk(CK), .q(g262), .d(g6042) );
  dff_311 DFF_223 ( .clk(CK), .q(g1840), .d(g8384) );
  dff_310 DFF_224 ( .clk(CK), .q(g70), .d(g6653) );
  dff_309 DFF_225 ( .clk(CK), .q(g318), .d(g257) );
  dff_308 DFF_226 ( .clk(CK), .q(g1356), .d(g5763) );
  dff_307 DFF_227 ( .clk(CK), .q(g794), .d(g5849) );
  dff_306 DFF_228 ( .clk(CK), .q(g36), .d(g10722) );
  dff_305 DFF_229 ( .clk(CK), .q(g302), .d(g6929) );
  dff_304 DFF_230 ( .clk(CK), .q(g342), .d(g11488) );
  dff_303 DFF_231 ( .clk(CK), .q(g1250), .d(g7299) );
  dff_302 DFF_232 ( .clk(CK), .q(g1163), .d(g4330) );
  dff_301 DFF_233 ( .clk(CK), .q(g1810), .d(g1958) );
  dff_300 DFF_234 ( .clk(CK), .q(g1032), .d(g7257) );
  dff_299 DFF_235 ( .clk(CK), .q(g1432), .d(g8775) );
  dff_298 DFF_236 ( .clk(CK), .q(g1053), .d(g7225) );
  dff_297 DFF_237 ( .clk(CK), .q(g1453), .d(g5770) );
  dff_296 DFF_238 ( .clk(CK), .q(g363), .d(g11486) );
  dff_295 DFF_239 ( .clk(CK), .q(g330), .d(g261) );
  dff_294 DFF_240 ( .clk(CK), .q(g1157), .d(g4338) );
  dff_293 DFF_241 ( .clk(CK), .q(g1357), .d(g4500) );
  dff_292 DFF_242 ( .clk(CK), .q(g35), .d(g10721) );
  dff_291 DFF_243 ( .clk(CK), .q(g928), .d(g8147) );
  dff_290 DFF_244 ( .clk(CK), .q(g261), .d(g6038) );
  dff_289 DFF_245 ( .clk(CK), .q(g516), .d(g11337) );
  dff_288 DFF_246 ( .clk(CK), .q(g254), .d(g6045) );
  dff_287 DFF_247 ( .clk(CK), .q(g778), .d(g7191) );
  dff_286 DFF_248 ( .clk(CK), .q(g861), .d(g826) );
  dff_285 DFF_249 ( .clk(CK), .q(g1627), .d(g8774) );
  dff_284 DFF_250 ( .clk(CK), .q(g1292), .d(g7293) );
  dff_283 DFF_251 ( .clk(CK), .q(g290), .d(g6907) );
  dff_282 DFF_252 ( .clk(CK), .q(g1850), .d(g4903) );
  dff_281 DFF_253 ( .clk(CK), .q(g770), .d(g6123) );
  dff_280 DFF_254 ( .clk(CK), .q(g1583), .d(g6506) );
  dff_279 DFF_255 ( .clk(CK), .q(g466), .d(g11376) );
  dff_278 DFF_256 ( .clk(CK), .q(g1561), .d(g6542) );
  dff_277 DFF_257 ( .clk(CK), .q(g1527), .d(g2807) );
  dff_276 DFF_258 ( .clk(CK), .q(g1546), .d(g6551) );
  dff_275 DFF_259 ( .clk(CK), .q(g287), .d(g6901) );
  dff_274 DFF_260 ( .clk(CK), .q(g560), .d(g10797) );
  dff_273 DFF_261 ( .clk(CK), .q(g617), .d(g8505) );
  dff_272 DFF_262 ( .clk(CK), .q(g17), .d(g4117) );
  dff_271 DFF_263 ( .clk(CK), .q(g336), .d(g11647) );
  dff_270 DFF_264 ( .clk(CK), .q(g456), .d(g11340) );
  dff_269 DFF_265 ( .clk(CK), .q(g305), .d(g253) );
  dff_268 DFF_266 ( .clk(CK), .q(g345), .d(g11625) );
  dff_267 DFF_267 ( .clk(CK), .q(g8), .d(g636) );
  dff_266 DFF_268 ( .clk(CK), .q(g1771), .d(g6502) );
  dff_265 DFF_269 ( .clk(CK), .q(g865), .d(n1272) );
  dff_264 DFF_270 ( .clk(CK), .q(g255), .d(g6049) );
  dff_263 DFF_271 ( .clk(CK), .q(g1945), .d(g8945) );
  dff_262 DFF_272 ( .clk(CK), .q(g1738), .d(g4231) );
  dff_261 DFF_273 ( .clk(CK), .q(g1478), .d(g8040) );
  dff_260 DFF_274 ( .clk(CK), .q(g1035), .d(g7203) );
  dff_259 DFF_275 ( .clk(CK), .q(g1959), .d(n1302) );
  dff_258 DFF_276 ( .clk(CK), .q(g1690), .d(g6155) );
  dff_257 DFF_277 ( .clk(CK), .q(g1482), .d(g8043) );
  dff_256 DFF_278 ( .clk(CK), .q(g1110), .d(g5173) );
  dff_255 DFF_279 ( .clk(CK), .q(g296), .d(g6916) );
  dff_254 DFF_280 ( .clk(CK), .q(g1663), .d(g10861) );
  dff_253 DFF_281 ( .clk(CK), .q(g700), .d(g8431) );
  dff_252 DFF_282 ( .clk(CK), .q(g1762), .d(g4309) );
  dff_251 DFF_283 ( .clk(CK), .q(g360), .d(g11485) );
  dff_250 DFF_284 ( .clk(CK), .q(g192), .d(g6334) );
  dff_249 DFF_285 ( .clk(CK), .q(g1657), .d(g10767) );
  dff_248 DFF_286 ( .clk(CK), .q(g722), .d(g8923) );
  dff_247 DFF_287 ( .clk(CK), .q(g61), .d(g7189) );
  dff_246 DFF_288 ( .clk(CK), .q(g566), .d(g10799) );
  dff_245 DFF_289 ( .clk(CK), .q(g1394), .d(g6747) );
  dff_244 DFF_290 ( .clk(CK), .q(g1089), .d(g6080) );
  dff_243 DFF_291 ( .clk(CK), .q(g883), .d(g3381) );
  dff_242 DFF_292 ( .clk(CK), .q(g1071), .d(g5910) );
  dff_241 DFF_293 ( .clk(CK), .q(g986), .d(g11393) );
  dff_240 DFF_294 ( .clk(CK), .q(g971), .d(g11349) );
  dff_239 DFF_295 ( .clk(CK), .q(g1955), .d(g83) );
  dff_238 DFF_296 ( .clk(CK), .q(g143), .d(g6439) );
  dff_237 DFF_297 ( .clk(CK), .q(g1814), .d(g9266) );
  dff_236 DFF_298 ( .clk(CK), .q(g1038), .d(g7245) );
  dff_235 DFF_299 ( .clk(CK), .q(g1212), .d(g1217) );
  dff_234 DFF_300 ( .clk(CK), .q(g1918), .d(g8940) );
  dff_233 DFF_301 ( .clk(CK), .q(g782), .d(g7705) );
  dff_232 DFF_302 ( .clk(CK), .q(g1822), .d(g9269) );
  dff_231 DFF_303 ( .clk(CK), .q(g237), .d(g6820) );
  dff_230 DFF_304 ( .clk(CK), .q(g746), .d(g756) );
  dff_229 DFF_305 ( .clk(CK), .q(g1062), .d(g7240) );
  dff_228 DFF_306 ( .clk(CK), .q(g1462), .d(g8042) );
  dff_227 DFF_307 ( .clk(CK), .q(g178), .d(g6759) );
  dff_226 DFF_308 ( .clk(CK), .q(g366), .d(g11487) );
  dff_225 DFF_309 ( .clk(CK), .q(g837), .d(g802) );
  dff_224 DFF_310 ( .clk(CK), .q(g599), .d(g9124) );
  dff_223 DFF_311 ( .clk(CK), .q(g1854), .d(g11293) );
  dff_222 DFF_312 ( .clk(CK), .q(g944), .d(g11298) );
  dff_221 DFF_313 ( .clk(CK), .q(g1941), .d(g8287) );
  dff_220 DFF_314 ( .clk(CK), .q(g170), .d(g8047) );
  dff_219 DFF_315 ( .clk(CK), .q(g1520), .d(g6205) );
  dff_218 DFF_316 ( .clk(CK), .q(g686), .d(g8885) );
  dff_217 DFF_317 ( .clk(CK), .q(g953), .d(g11305) );
  dff_216 DFF_318 ( .clk(CK), .q(g1958), .d(g5556) );
  dff_215 DFF_319 ( .clk(CK), .q(g40), .d(g10664) );
  dff_214 DFF_320 ( .clk(CK), .q(g1765), .d(g2478) );
  dff_213 DFF_321 ( .clk(CK), .q(g1733), .d(g10711) );
  dff_212 DFF_322 ( .clk(CK), .q(g1270), .d(g7303) );
  dff_211 DFF_323 ( .clk(CK), .q(g1610), .d(g5194) );
  dff_210 DFF_324 ( .clk(CK), .q(g1796), .d(g7541) );
  dff_209 DFF_325 ( .clk(CK), .q(g1324), .d(g11607) );
  dff_208 DFF_326 ( .clk(CK), .q(g1540), .d(g6541) );
  dff_207 DFF_327 ( .clk(CK), .q(g1377), .d(g6827) );
  dff_206 DFF_328 ( .clk(CK), .q(g1206), .d(g4114) );
  dff_205 DFF_329 ( .clk(CK), .q(g491), .d(g11332) );
  dff_204 DFF_330 ( .clk(CK), .q(g1849), .d(g4902) );
  dff_203 DFF_331 ( .clk(CK), .q(g213), .d(g6828) );
  dff_202 DFF_332 ( .clk(CK), .q(g1781), .d(g6516) );
  dff_201 DFF_333 ( .clk(CK), .q(g1900), .d(g8938) );
  dff_200 DFF_334 ( .clk(CK), .q(g1245), .d(g7298) );
  dff_199 DFF_335 ( .clk(CK), .q(g108), .d(g11561) );
  dff_198 DFF_336 ( .clk(CK), .q(g630), .d(g6672) );
  dff_197 DFF_337 ( .clk(CK), .q(g148), .d(g8048) );
  dff_196 DFF_338 ( .clk(CK), .q(g833), .d(g798) );
  dff_195 DFF_339 ( .clk(CK), .q(g1923), .d(g8285) );
  dff_194 DFF_340 ( .clk(CK), .q(g936), .d(g8254) );
  dff_193 DFF_341 ( .clk(CK), .q(g1215), .d(g5229) );
  dff_192 DFF_342 ( .clk(CK), .q(g1314), .d(g11604) );
  dff_191 DFF_343 ( .clk(CK), .q(g849), .d(g814) );
  dff_190 DFF_344 ( .clk(CK), .q(g1336), .d(g11636) );
  dff_189 DFF_345 ( .clk(CK), .q(g272), .d(g6910) );
  dff_188 DFF_346 ( .clk(CK), .q(g1806), .d(g8173) );
  dff_187 DFF_347 ( .clk(CK), .q(g826), .d(g8245) );
  dff_186 DFF_348 ( .clk(CK), .q(g1065), .d(g7242) );
  dff_185 DFF_349 ( .clk(CK), .q(g1887), .d(g8281) );
  dff_184 DFF_350 ( .clk(CK), .q(g37), .d(g10724) );
  dff_183 DFF_351 ( .clk(CK), .q(g968), .d(g11314) );
  dff_182 DFF_352 ( .clk(CK), .q(g1845), .d(g4905) );
  dff_181 DFF_353 ( .clk(CK), .q(g1137), .d(g4484) );
  dff_180 DFF_354 ( .clk(CK), .q(g1891), .d(g8937) );
  dff_179 DFF_355 ( .clk(CK), .q(g1255), .d(g7300) );
  dff_178 DFF_356 ( .clk(CK), .q(g257), .d(g6002) );
  dff_177 DFF_357 ( .clk(CK), .q(g874), .d(n1186) );
  dff_176 DFF_358 ( .clk(CK), .q(g591), .d(g9110) );
  dff_175 DFF_359 ( .clk(CK), .q(g731), .d(g8926) );
  dff_174 DFF_360 ( .clk(CK), .q(g636), .d(g8631) );
  dff_173 DFF_361 ( .clk(CK), .q(g1218), .d(g7632) );
  dff_172 DFF_362 ( .clk(CK), .q(g605), .d(g9150) );
  dff_171 DFF_363 ( .clk(CK), .q(g79), .d(g6531) );
  dff_170 DFF_364 ( .clk(CK), .q(g182), .d(g6786) );
  dff_169 DFF_365 ( .clk(CK), .q(g950), .d(g11303) );
  dff_168 DFF_366 ( .clk(CK), .q(g1129), .d(g4477) );
  dff_167 DFF_367 ( .clk(CK), .q(g857), .d(g822) );
  dff_166 DFF_368 ( .clk(CK), .q(g448), .d(g11258) );
  dff_165 DFF_369 ( .clk(CK), .q(g1828), .d(g9272) );
  dff_164 DFF_370 ( .clk(CK), .q(g1727), .d(g10773) );
  dff_163 DFF_371 ( .clk(CK), .q(g1592), .d(g6470) );
  dff_162 DFF_372 ( .clk(CK), .q(g1703), .d(g5083) );
  dff_161 DFF_373 ( .clk(CK), .q(g1932), .d(g8286) );
  dff_160 DFF_374 ( .clk(CK), .q(g1624), .d(g8773) );
  dff_159 DFF_375 ( .clk(CK), .q(g26), .d(n1256) );
  dff_158 DFF_376 ( .clk(CK), .q(g1068), .d(g6054) );
  dff_157 DFF_377 ( .clk(CK), .q(g578), .d(g101) );
  dff_156 DFF_378 ( .clk(CK), .q(g440), .d(g11260) );
  dff_155 DFF_379 ( .clk(CK), .q(g476), .d(g11338) );
  dff_154 DFF_380 ( .clk(CK), .q(g119), .d(g5918) );
  dff_153 DFF_381 ( .clk(CK), .q(g668), .d(g8922) );
  dff_152 DFF_382 ( .clk(CK), .q(g139), .d(g8049) );
  dff_151 DFF_383 ( .clk(CK), .q(g1149), .d(g4342) );
  dff_150 DFF_384 ( .clk(CK), .q(g34), .d(g10720) );
  dff_149 DFF_385 ( .clk(CK), .q(g1848), .d(g6755) );
  dff_148 DFF_386 ( .clk(CK), .q(g263), .d(g6897) );
  dff_147 DFF_387 ( .clk(CK), .q(g818), .d(g7709) );
  dff_146 DFF_388 ( .clk(CK), .q(g1747), .d(g4255) );
  dff_145 DFF_389 ( .clk(CK), .q(g802), .d(g5543) );
  dff_144 DFF_390 ( .clk(CK), .q(g275), .d(g6915) );
  dff_143 DFF_391 ( .clk(CK), .q(g1524), .d(g6513) );
  dff_142 DFF_392 ( .clk(CK), .q(g1577), .d(g6480) );
  dff_141 DFF_393 ( .clk(CK), .q(g810), .d(g6733) );
  dff_140 DFF_394 ( .clk(CK), .q(g391), .d(g11264) );
  dff_139 DFF_395 ( .clk(CK), .q(g658), .d(g8973) );
  dff_138 DFF_396 ( .clk(CK), .q(g1386), .d(g6833) );
  dff_137 DFF_397 ( .clk(CK), .q(g253), .d(g5996) );
  dff_136 DFF_398 ( .clk(CK), .q(g875), .d(n1175) );
  dff_135 DFF_399 ( .clk(CK), .q(g1125), .d(g4473) );
  dff_134 DFF_400 ( .clk(CK), .q(g201), .d(g5755) );
  dff_133 DFF_401 ( .clk(CK), .q(g1280), .d(g7295) );
  dff_132 DFF_402 ( .clk(CK), .q(g1083), .d(g6068) );
  dff_131 DFF_403 ( .clk(CK), .q(g650), .d(g7137) );
  dff_130 DFF_404 ( .clk(CK), .q(g1636), .d(g8779) );
  dff_129 DFF_405 ( .clk(CK), .q(g853), .d(g818) );
  dff_128 DFF_406 ( .clk(CK), .q(g421), .d(g11270) );
  dff_127 DFF_407 ( .clk(CK), .q(g762), .d(g5529) );
  dff_126 DFF_408 ( .clk(CK), .q(g956), .d(g11306) );
  dff_125 DFF_409 ( .clk(CK), .q(g378), .d(g11291) );
  dff_124 DFF_410 ( .clk(CK), .q(g1756), .d(g4283) );
  dff_123 DFF_411 ( .clk(CK), .q(g589), .d(g29) );
  dff_122 DFF_412 ( .clk(CK), .q(g841), .d(g806) );
  dff_121 DFF_413 ( .clk(CK), .q(g1027), .d(g6894) );
  dff_120 DFF_414 ( .clk(CK), .q(g1003), .d(g6902) );
  dff_119 DFF_415 ( .clk(CK), .q(g1403), .d(g8765) );
  dff_118 DFF_416 ( .clk(CK), .q(g1145), .d(g4498) );
  dff_117 DFF_417 ( .clk(CK), .q(g1107), .d(g5148) );
  dff_116 DFF_418 ( .clk(CK), .q(g1223), .d(g7581) );
  dff_115 DFF_419 ( .clk(CK), .q(g406), .d(g11267) );
  dff_114 DFF_420 ( .clk(CK), .q(g1811), .d(g10936) );
  dff_113 DFF_421 ( .clk(CK), .q(g1642), .d(g10784) );
  dff_112 DFF_422 ( .clk(CK), .q(g1047), .d(g7211) );
  dff_111 DFF_423 ( .clk(CK), .q(g1654), .d(g10765) );
  dff_110 DFF_424 ( .clk(CK), .q(g197), .d(g6332) );
  dff_109 DFF_425 ( .clk(CK), .q(g1595), .d(g6479) );
  dff_108 DFF_426 ( .clk(CK), .q(g1537), .d(g6537) );
  dff_107 DFF_427 ( .clk(CK), .q(g727), .d(g8434) );
  dff_106 DFF_428 ( .clk(CK), .q(g999), .d(g6908) );
  dff_105 DFF_429 ( .clk(CK), .q(g798), .d(g6243) );
  dff_104 DFF_430 ( .clk(CK), .q(g481), .d(g11324) );
  dff_103 DFF_431 ( .clk(CK), .q(g754), .d(g3462) );
  dff_102 DFF_432 ( .clk(CK), .q(g1330), .d(g11609) );
  dff_101 DFF_433 ( .clk(CK), .q(g845), .d(g810) );
  dff_100 DFF_434 ( .clk(CK), .q(g790), .d(g8244) );
  dff_99 DFF_435 ( .clk(CK), .q(g1512), .d(g8194) );
  dff_98 DFF_436 ( .clk(CK), .q(g114), .d(g113) );
  dff_97 DFF_437 ( .clk(CK), .q(g1490), .d(g8052) );
  dff_96 DFF_438 ( .clk(CK), .q(g1166), .d(g4325) );
  dff_95 DFF_439 ( .clk(CK), .q(g1056), .d(g7231) );
  dff_94 DFF_440 ( .clk(CK), .q(g348), .d(g11481) );
  dff_93 DFF_441 ( .clk(CK), .q(g868), .d(g874) );
  dff_92 DFF_442 ( .clk(CK), .q(g1260), .d(g7301) );
  dff_91 DFF_443 ( .clk(CK), .q(g260), .d(g6035) );
  dff_90 DFF_444 ( .clk(CK), .q(g131), .d(g8059) );
  dff_89 DFF_445 ( .clk(CK), .q(g7), .d(g1854) );
  dff_88 DFF_446 ( .clk(CK), .q(g258), .d(g6015) );
  dff_87 DFF_447 ( .clk(CK), .q(g521), .d(g11330) );
  dff_86 DFF_448 ( .clk(CK), .q(g1318), .d(g11605) );
  dff_85 DFF_449 ( .clk(CK), .q(g1872), .d(g8921) );
  dff_84 DFF_450 ( .clk(CK), .q(g677), .d(g8883) );
  dff_83 DFF_451 ( .clk(CK), .q(g582), .d(g28) );
  dff_82 DFF_452 ( .clk(CK), .q(g1393), .d(g6163) );
  dff_81 DFF_453 ( .clk(CK), .q(g1549), .d(g6523) );
  dff_80 DFF_454 ( .clk(CK), .q(g947), .d(g11300) );
  dff_79 DFF_455 ( .clk(CK), .q(g1834), .d(g9555) );
  dff_78 DFF_456 ( .clk(CK), .q(g1598), .d(g6481) );
  dff_77 DFF_457 ( .clk(CK), .q(g1121), .d(g4471) );
  dff_76 DFF_458 ( .clk(CK), .q(g1321), .d(g11606) );
  dff_75 DFF_459 ( .clk(CK), .q(g506), .d(g11335) );
  dff_74 DFF_460 ( .clk(CK), .q(g546), .d(g10791) );
  dff_73 DFF_461 ( .clk(CK), .q(g1909), .d(g8939) );
  dff_72 DFF_462 ( .clk(CK), .q(g755), .d(g83) );
  dff_71 DFF_463 ( .clk(CK), .q(g1552), .d(g6529) );
  dff_70 DFF_464 ( .clk(CK), .q(g584), .d(g101) );
  dff_69 DFF_465 ( .clk(CK), .q(g1687), .d(g10776) );
  dff_68 DFF_466 ( .clk(CK), .q(g1586), .d(g6514) );
  dff_67 DFF_467 ( .clk(CK), .q(g324), .d(g259) );
  dff_66 DFF_468 ( .clk(CK), .q(g1141), .d(g4490) );
  dff_65 DFF_469 ( .clk(CK), .q(g1570), .d(g2807) );
  dff_64 DFF_470 ( .clk(CK), .q(g1341), .d(g11639) );
  dff_63 DFF_471 ( .clk(CK), .q(g1710), .d(g4089) );
  dff_62 DFF_472 ( .clk(CK), .q(g1645), .d(g10785) );
  dff_61 DFF_473 ( .clk(CK), .q(g115), .d(g6179) );
  dff_60 DFF_474 ( .clk(CK), .q(g135), .d(g8053) );
  dff_59 DFF_475 ( .clk(CK), .q(g525), .d(g11329) );
  dff_58 DFF_476 ( .clk(CK), .q(g581), .d(g104) );
  dff_57 DFF_477 ( .clk(CK), .q(g1607), .d(g6515) );
  dff_56 DFF_478 ( .clk(CK), .q(g321), .d(g258) );
  dff_55 DFF_479 ( .clk(CK), .q(g67), .d(g7204) );
  dff_54 DFF_480 ( .clk(CK), .q(g1275), .d(g11443) );
  dff_53 DFF_481 ( .clk(CK), .q(g1311), .d(g11603) );
  dff_52 DFF_482 ( .clk(CK), .q(g1615), .d(g8770) );
  dff_51 DFF_483 ( .clk(CK), .q(g382), .d(g11292) );
  dff_50 DFF_484 ( .clk(CK), .q(g1374), .d(g6331) );
  dff_49 DFF_485 ( .clk(CK), .q(g266), .d(g6900) );
  dff_48 DFF_486 ( .clk(CK), .q(g1284), .d(g7294) );
  dff_47 DFF_487 ( .clk(CK), .q(g1380), .d(g6829) );
  dff_46 DFF_488 ( .clk(CK), .q(g673), .d(g8428) );
  dff_45 DFF_489 ( .clk(CK), .q(g1853), .d(g4904) );
  dff_44 DFF_490 ( .clk(CK), .q(g162), .d(g8054) );
  dff_43 DFF_491 ( .clk(CK), .q(g411), .d(g11268) );
  dff_42 DFF_492 ( .clk(CK), .q(g431), .d(g11262) );
  dff_41 DFF_493 ( .clk(CK), .q(g1905), .d(g8283) );
  dff_40 DFF_494 ( .clk(CK), .q(g1515), .d(g6193) );
  dff_39 DFF_495 ( .clk(CK), .q(g1630), .d(g8776) );
  dff_38 DFF_496 ( .clk(CK), .q(g49), .d(g7143) );
  dff_37 DFF_497 ( .clk(CK), .q(g991), .d(g6898) );
  dff_36 DFF_498 ( .clk(CK), .q(g1300), .d(g7291) );
  dff_35 DFF_499 ( .clk(CK), .q(g339), .d(g11478) );
  dff_34 DFF_500 ( .clk(CK), .q(g256), .d(g6000) );
  dff_33 DFF_501 ( .clk(CK), .q(g1750), .d(g4264) );
  dff_32 DFF_502 ( .clk(CK), .q(g585), .d(g102) );
  dff_31 DFF_503 ( .clk(CK), .q(g1440), .d(g8768) );
  dff_30 DFF_504 ( .clk(CK), .q(g1666), .d(g10863) );
  dff_29 DFF_505 ( .clk(CK), .q(g1528), .d(g6522) );
  dff_28 DFF_506 ( .clk(CK), .q(g1351), .d(g11641) );
  dff_27 DFF_507 ( .clk(CK), .q(g1648), .d(g10780) );
  dff_26 DFF_508 ( .clk(CK), .q(g127), .d(g8044) );
  dff_25 DFF_509 ( .clk(CK), .q(g1618), .d(g11579) );
  dff_24 DFF_510 ( .clk(CK), .q(g1235), .d(g7296) );
  dff_23 DFF_511 ( .clk(CK), .q(g299), .d(g6923) );
  dff_22 DFF_512 ( .clk(CK), .q(g435), .d(g11261) );
  dff_21 DFF_513 ( .clk(CK), .q(g64), .d(g6638) );
  dff_20 DFF_514 ( .clk(CK), .q(g1555), .d(g6534) );
  dff_19 DFF_515 ( .clk(CK), .q(g995), .d(g6895) );
  dff_18 DFF_516 ( .clk(CK), .q(g1621), .d(g8771) );
  dff_17 DFF_517 ( .clk(CK), .q(g1113), .d(g4506) );
  dff_16 DFF_518 ( .clk(CK), .q(g643), .d(g7441) );
  dff_15 DFF_519 ( .clk(CK), .q(g1494), .d(g8055) );
  dff_14 DFF_520 ( .clk(CK), .q(g1567), .d(g6468) );
  dff_13 DFF_521 ( .clk(CK), .q(g691), .d(g8430) );
  dff_12 DFF_522 ( .clk(CK), .q(g534), .d(g11327) );
  dff_11 DFF_523 ( .clk(CK), .q(g1776), .d(g6508) );
  dff_10 DFF_524 ( .clk(CK), .q(g569), .d(g10717) );
  dff_9 DFF_525 ( .clk(CK), .q(g1160), .d(g4334) );
  dff_8 DFF_526 ( .clk(CK), .q(g1360), .d(n1195) );
  dff_7 DFF_527 ( .clk(CK), .q(g1050), .d(g7218) );
  dff_6 DFF_528 ( .clk(CK), .q(g1), .d(g6679) );
  dff_5 DFF_529 ( .clk(CK), .q(g511), .d(g11336) );
  dff_4 DFF_530 ( .clk(CK), .q(g1724), .d(g10771) );
  dff_3 DFF_531 ( .clk(CK), .q(g12), .d(g5445) );
  dff_2 DFF_532 ( .clk(CK), .q(g1878), .d(g8559) );
  dff_1 DFF_533 ( .clk(CK), .q(g73), .d(g7219) );
  and2_0 AND2_0 ( .c(g11103), .b(g2250), .a(g10937) );
  and2_1553 AND2_1 ( .c(g9900), .b(g9088), .a(n1307) );
  and2_1552 AND2_2 ( .c(g11095), .b(g845), .a(g10950) );
  and2_1551 AND2_3 ( .c(g3880), .b(n1071), .a(n1097) );
  and2_1550 AND2_4 ( .c(g4973), .b(g1645), .a(n1202) );
  and2_1549 AND2_5 ( .c(g7389), .b(g5852), .a(g3880) );
  and2_1548 AND2_6 ( .c(g7888), .b(g7465), .a(n1253) );
  and2_1547 AND2_7 ( .c(g4969), .b(g1642), .a(n1202) );
  and2_1546 AND2_8 ( .c(g8224), .b(g1882), .a(n1210) );
  and2_1545 AND2_9 ( .c(g2892), .b(n1059), .a(n1157) );
  and2_1544 AND2_10 ( .c(g5686), .b(g158), .a(g5361) );
  and2_1543 AND2_11 ( .c(g10308), .b(g10013), .a(g8574) );
  and2_1542 AND2_12 ( .c(g4123), .b(n1339), .a(n1103) );
  and2_1541 AND2_13 ( .c(g8120), .b(g1909), .a(n1210) );
  and2_1540 AND2_14 ( .c(g6788), .b(g287), .a(n1221) );
  and2_1539 AND2_15 ( .c(g5598), .b(g778), .a(g4824) );
  and2_1538 AND2_16 ( .c(g9694), .b(g278), .a(n1171) );
  and2_1537 AND2_17 ( .c(g10495), .b(n1167), .a(n1071) );
  and2_1536 AND2_18 ( .c(g2945), .b(n1337), .a(g1684) );
  and2_1535 AND2_19 ( .c(g11190), .b(g4752), .a(n1350) );
  and2_1534 AND2_20 ( .c(g8789), .b(g8639), .a(n1213) );
  and2_1533 AND2_21 ( .c(g9852), .b(g9728), .a(g9563) );
  and2_1532 AND2_22 ( .c(g5625), .b(g1053), .a(n1368) );
  and2_1531 AND2_23 ( .c(g4875), .b(g995), .a(n1369) );
  and2_1530 AND2_24 ( .c(g9701), .b(g1574), .a(n1190) );
  and2_1529 AND2_25 ( .c(g7138), .b(g5201), .a(n1199) );
  and2_1528 AND2_26 ( .c(g10752), .b(g10599), .a(g3586) );
  and2_1527 AND2_27 ( .c(g11211), .b(g11058), .a(g3209) );
  and2_1526 AND2_28 ( .c(g11024), .b(g435), .a(n1346) );
  and2_1525 AND2_29 ( .c(g8547), .b(g8307), .a(g7246) );
  and2_1524 AND2_30 ( .c(g10669), .b(g10408), .a(n1224) );
  and2_1523 AND2_31 ( .c(g7707), .b(g691), .a(g6488) );
  and2_1522 AND2_32 ( .c(g4884), .b(g3813), .a(g1845) );
  and2_1521 AND2_33 ( .c(g4839), .b(g225), .a(n1386) );
  and2_1520 AND2_34 ( .c(g9870), .b(g1561), .a(g9324) );
  and2_1519 AND2_35 ( .c(g6640), .b(g86), .a(n1316) );
  and2_1518 AND2_36 ( .c(g9650), .b(g986), .a(n1330) );
  and2_1517 AND2_37 ( .c(g5687), .b(g139), .a(g5361) );
  and2_1516 AND2_38 ( .c(g7957), .b(g79), .a(n1383) );
  and2_1515 AND2_39 ( .c(g3512), .b(n1076), .a(g1845) );
  and2_1514 AND2_40 ( .c(g8244), .b(g7054), .a(n1286) );
  and2_1513 AND2_41 ( .c(g7449), .b(g6548), .a(n1264) );
  and2_1512 AND2_42 ( .c(g4235), .b(g1011), .a(n1372) );
  and2_1511 AND2_43 ( .c(g4343), .b(g345), .a(g3586) );
  and2_1510 AND2_44 ( .c(g11296), .b(g4561), .a(n1351) );
  and2_1509 AND2_45 ( .c(g9594), .b(g1), .a(n1331) );
  and2_1508 AND2_46 ( .c(g6829), .b(g213), .a(g5354) );
  and2_1507 AND2_47 ( .c(g4334), .b(g1160), .a(g109) );
  and2_1506 AND2_48 ( .c(g9943), .b(g9923), .a(n1320) );
  and2_1505 AND2_49 ( .c(g5525), .b(g1721), .a(n1185) );
  and2_1504 AND2_50 ( .c(g4548), .b(g440), .a(g109) );
  and3_0 AND3_0 ( .d(g8876), .c(n1252), .b(n1307), .a(n1281) );
  and2_1503 AND2_51 ( .c(g6733), .b(g4488), .a(n1277) );
  and2_1502 AND2_52 ( .c(g4804), .b(g476), .a(g109) );
  and2_1501 AND2_53 ( .c(g10705), .b(g10564), .a(n1367) );
  and2_1500 AND2_54 ( .c(g9934), .b(g9913), .a(g9624) );
  and2_1499 AND2_55 ( .c(g6225), .b(g566), .a(n1375) );
  and2_1498 AND2_56 ( .c(g6324), .b(g1240), .a(n1322) );
  and2_1497 AND2_57 ( .c(g10686), .b(g10385), .a(g3863) );
  and2_1496 AND2_58 ( .c(g6540), .b(g1223), .a(n1180) );
  and2_1495 AND2_59 ( .c(g8663), .b(g8270), .a(n1367) );
  and2_1494 AND2_60 ( .c(g11581), .b(g1308), .a(n1198) );
  and2_1493 AND2_61 ( .c(g6206), .b(g560), .a(n1370) );
  and2_1492 AND2_62 ( .c(g4518), .b(g452), .a(g109) );
  and2_1491 AND2_63 ( .c(g3989), .b(g248), .a(n1386) );
  and2_1490 AND2_64 ( .c(g7730), .b(g7260), .a(n1102) );
  and2_1489 AND2_65 ( .c(g5174), .b(g1235), .a(g109) );
  and2_1488 AND2_66 ( .c(g7504), .b(n1384), .a(g67) );
  and2_1487 AND2_67 ( .c(g7185), .b(g1887), .a(g6003) );
  and2_1486 AND2_68 ( .c(g2563), .b(I5689), .a(I5690) );
  and2_1485 AND2_69 ( .c(g7881), .b(g5295), .a(n1388) );
  and2_1484 AND2_70 ( .c(g11070), .b(n1107), .a(g10788) );
  and2_1483 AND2_71 ( .c(g9859), .b(g9736), .a(g9573) );
  and3_48 AND3_1 ( .d(g8877), .c(n1249), .b(n1307), .a(n1281) );
  and2_1482 AND2_72 ( .c(g11590), .b(g2274), .a(g11561) );
  and2_1481 AND2_73 ( .c(g6199), .b(g557), .a(n1370) );
  and2_1480 AND2_74 ( .c(g9266), .b(g8932), .a(n1386) );
  and2_1479 AND2_75 ( .c(g5545), .b(g1730), .a(n1185) );
  and2_1478 AND2_76 ( .c(g5180), .b(g814), .a(g810) );
  and2_1477 AND2_77 ( .c(g5591), .b(g1615), .a(n1390) );
  and2_1476 AND2_78 ( .c(g8556), .b(g8412), .a(g7638) );
  and2_1475 AND2_79 ( .c(g11094), .b(g374), .a(n1163) );
  and2_1474 AND2_80 ( .c(g5853), .b(g5044), .a(g1927) );
  and2_1473 AND2_81 ( .c(g6245), .b(g575), .a(n1370) );
  and2_1472 AND2_82 ( .c(g4360), .b(g1861), .a(n1124) );
  and3_47 AND3_2 ( .d(g8930), .c(n1290), .b(n1307), .a(n1266) );
  and2_1471 AND2_83 ( .c(g5507), .b(g563), .a(n1391) );
  and2_1470 AND2_84 ( .c(g11150), .b(g3087), .a(g10788) );
  and2_1469 AND2_85 ( .c(g8464), .b(g8302), .a(g7246) );
  and2_1468 AND2_86 ( .c(g9692), .b(g272), .a(n1171) );
  and2_1467 AND2_87 ( .c(g4996), .b(g1428), .a(g4682) );
  and2_1466 AND2_88 ( .c(g7131), .b(g5174), .a(n1199) );
  and2_1465 AND2_89 ( .c(g11019), .b(g421), .a(n1346) );
  and2_1464 AND2_90 ( .c(g9960), .b(g9951), .a(n1319) );
  and2_1463 AND2_91 ( .c(g11196), .b(g4770), .a(n1352) );
  and2_1462 AND2_92 ( .c(g11018), .b(g6485), .a(n1346) );
  and2_1461 AND2_93 ( .c(g6819), .b(g243), .a(g5354) );
  and2_1460 AND2_94 ( .c(g10595), .b(g10550), .a(n1159) );
  and2_1459 AND2_95 ( .c(g10494), .b(g10433), .a(n1071) );
  and2_1458 AND2_96 ( .c(g10623), .b(g10544), .a(n1159) );
  and2_1457 AND2_97 ( .c(g4878), .b(g1868), .a(n1124) );
  and2_1456 AND2_98 ( .c(g5204), .b(g4838), .a(n1158) );
  and2_1455 AND2_99 ( .c(g8844), .b(g8609), .a(n1233) );
  and2_1454 AND2_100 ( .c(g6701), .b(g6185), .a(n1367) );
  and2_1453 AND2_101 ( .c(g10782), .b(g10725), .a(n1202) );
  and2_1452 AND2_102 ( .c(g5100), .b(g1791), .a(n1202) );
  and2_1451 AND2_103 ( .c(g4882), .b(g1089), .a(n1367) );
  and2_1450 AND2_104 ( .c(g8731), .b(g8236), .a(n1384) );
  and2_1449 AND2_105 ( .c(g6215), .b(g1504), .a(g5128) );
  and2_1448 AND2_106 ( .c(g6886), .b(g1932), .a(g6003) );
  and2_1447 AND2_107 ( .c(g3586), .b(g1703), .a(n1301) );
  and2_1446 AND2_108 ( .c(g8557), .b(g8415), .a(g7638) );
  and3_46 AND3_3 ( .d(g8966), .c(n1284), .b(n1307), .a(n1274) );
  and2_1445 AND2_109 ( .c(g8071), .b(g691), .a(n1251) );
  and2_1444 AND2_110 ( .c(g11597), .b(g11549), .a(g4421) );
  and2_1443 AND2_111 ( .c(g9828), .b(g9722), .a(g9785) );
  and2_1442 AND2_112 ( .c(g2918), .b(n1337), .a(g1672) );
  and2_1441 AND2_113 ( .c(g9830), .b(g9725), .a(g9785) );
  and3_45 AND3_4 ( .d(g8955), .c(n1283), .b(n1307), .a(n1266) );
  and2_1440 AND2_114 ( .c(g9592), .b(g4), .a(n1331) );
  and2_1439 AND2_115 ( .c(g5123), .b(g1618), .a(n1370) );
  and2_1438 AND2_116 ( .c(g7059), .b(g6078), .a(n1236) );
  and2_1437 AND2_117 ( .c(g8254), .b(g936), .a(n1209) );
  and2_1436 AND2_118 ( .c(g7459), .b(n1384), .a(g55) );
  and2_1435 AND2_119 ( .c(g11102), .b(g861), .a(g10950) );
  and2_1434 AND2_120 ( .c(g7718), .b(g709), .a(g6488) );
  and2_1433 AND2_121 ( .c(g7535), .b(n1384), .a(g49) );
  and2_1432 AND2_122 ( .c(g9703), .b(g1577), .a(n1190) );
  and2_1431 AND2_123 ( .c(g5528), .b(g569), .a(n1391) );
  and2_1430 AND2_124 ( .c(g5151), .b(n1295), .a(g109) );
  and2_1429 AND2_125 ( .c(g9932), .b(g9911), .a(g9624) );
  and2_1428 AND2_126 ( .c(g5530), .b(g1636), .a(n1371) );
  and2_1427 AND2_127 ( .c(g3506), .b(g986), .a(g2760) );
  and2_1426 AND2_128 ( .c(g8769), .b(g8629), .a(g5151) );
  and2_1425 AND2_129 ( .c(g6887), .b(g6187), .a(n1267) );
  and2_1424 AND2_130 ( .c(g6228), .b(g5605), .a(g713) );
  and2_1423 AND2_131 ( .c(g6322), .b(g1275), .a(n1322) );
  and2_1422 AND2_132 ( .c(g3111), .b(I6337), .a(I6338) );
  and3_44 AND3_5 ( .d(g8967), .c(n1271), .b(n1307), .a(n1274) );
  and2_1421 AND2_133 ( .c(g5010), .b(g1458), .a(g4640) );
  and2_1420 AND2_134 ( .c(g3275), .b(g115), .a(n1386) );
  and2_1419 AND2_135 ( .c(g10809), .b(n1196), .a(n1346) );
  and2_1418 AND2_136 ( .c(g2895), .b(n1337), .a(g1678) );
  and2_1417 AND2_137 ( .c(g7721), .b(g736), .a(g6488) );
  and2_1416 AND2_138 ( .c(g9866), .b(g1549), .a(g9324) );
  and2_1415 AND2_139 ( .c(g9716), .b(g1534), .a(n1207) );
  and2_1414 AND2_140 ( .c(g10808), .b(g10744), .a(g3829) );
  and2_1413 AND2_141 ( .c(g3374), .b(g1231), .a(g3047) );
  and2_1412 AND2_142 ( .c(g4492), .b(g1786), .a(g3685) );
  and2_1411 AND2_143 ( .c(g8822), .b(g8614), .a(n1233) );
  and2_1410 AND2_144 ( .c(g10560), .b(g10369), .a(n1159) );
  and3_43 AND3_6 ( .d(g11456), .c(n1228), .b(n1287), .a(n1275) );
  and2_1409 AND2_145 ( .c(g9848), .b(g9724), .a(g9557) );
  and2_1408 AND2_146 ( .c(g4714), .b(g646), .a(n1089) );
  and2_1407 AND2_147 ( .c(g6550), .b(g1231), .a(n1180) );
  and2_1406 AND2_148 ( .c(g5172), .b(g822), .a(g818) );
  and2_1405 AND2_149 ( .c(g10642), .b(g10385), .a(g3829) );
  and2_1404 AND2_150 ( .c(g3284), .b(g2531), .a(g677) );
  and2_1403 AND2_151 ( .c(g9699), .b(g284), .a(n1171) );
  and2_1402 AND2_152 ( .c(g9855), .b(g302), .a(g9313) );
  and2_1401 AND2_153 ( .c(g5618), .b(g1630), .a(n1391) );
  and2_1400 AND2_154 ( .c(g6891), .b(g1950), .a(g6003) );
  and2_1399 AND2_155 ( .c(g7940), .b(g5319), .a(n1367) );
  and2_1398 AND2_156 ( .c(g11085), .b(g312), .a(n1352) );
  and2_1397 AND2_157 ( .c(g4736), .b(g396), .a(g109) );
  and2_1396 AND2_158 ( .c(g4968), .b(g1432), .a(g4682) );
  and2_1395 AND2_159 ( .c(g8837), .b(g8646), .a(n1213) );
  and2_1394 AND2_160 ( .c(g9644), .b(g1182), .a(g9125) );
  and2_1393 AND2_161 ( .c(g5804), .b(g1546), .a(n1229) );
  and2_1392 AND2_162 ( .c(g8462), .b(g8300), .a(g7246) );
  and4_0 AND4_0 ( .e(I6330), .d(n1138), .c(n1068), .b(n1087), .a(n1046) );
  and2_1391 AND2_163 ( .c(g11156), .b(g333), .a(n1352) );
  and2_1390 AND2_164 ( .c(g6342), .b(g293), .a(n1221) );
  and2_1389 AND2_165 ( .c(g9867), .b(g1552), .a(g9324) );
  and2_1388 AND2_166 ( .c(g9717), .b(g1537), .a(n1207) );
  and2_1387 AND2_167 ( .c(g4871), .b(g1864), .a(n1124) );
  and2_1386 AND2_168 ( .c(g10454), .b(g10435), .a(n1071) );
  and2_1385 AND2_169 ( .c(g4722), .b(g426), .a(g109) );
  and2_1384 AND2_170 ( .c(g7741), .b(g5824), .a(g3880) );
  and2_1383 AND2_171 ( .c(g4500), .b(g1357), .a(n1371) );
  and2_1382 AND2_172 ( .c(g9386), .b(g1327), .a(n1325) );
  and2_1381 AND2_173 ( .c(g8842), .b(g8607), .a(n1233) );
  and2_1380 AND2_174 ( .c(g9599), .b(g8), .a(n1331) );
  and2_1379 AND2_175 ( .c(g9274), .b(g8974), .a(g48) );
  and2_1378 AND2_176 ( .c(g5518), .b(g566), .a(n1391) );
  and2_1377 AND2_177 ( .c(g9614), .b(g1197), .a(g9111) );
  and2_1376 AND2_178 ( .c(g4838), .b(g3275), .a(g4122) );
  and2_1375 AND2_179 ( .c(g9125), .b(g8966), .a(g48) );
  and2_1374 AND2_180 ( .c(g7217), .b(g4610), .a(n1276) );
  and2_1373 AND2_181 ( .c(g11557), .b(g1791), .a(g11519) );
  and2_1372 AND2_182 ( .c(g2911), .b(n1337), .a(g1675) );
  and2_1371 AND2_183 ( .c(g11210), .b(g10886), .a(n1254) );
  and2_1370 AND2_184 ( .c(g7466), .b(n1384), .a(g58) );
  and2_1369 AND2_185 ( .c(g9939), .b(g9918), .a(n1320) );
  and2_1368 AND2_186 ( .c(g11279), .b(g4784), .a(n1352) );
  and3_42 AND3_7 ( .d(g10518), .c(g10513), .b(g10440), .a(I16145) );
  and2_1367 AND2_187 ( .c(g4477), .b(g1129), .a(g109) );
  and2_1366 AND2_188 ( .c(g8708), .b(n1234), .a(g8488) );
  and2_1365 AND2_189 ( .c(g7055), .b(g5004), .a(n1199) );
  and2_1364 AND2_190 ( .c(g5264), .b(g1095), .a(n1161) );
  and2_1363 AND2_191 ( .c(g6329), .b(g1265), .a(n1322) );
  and2_1362 AND2_192 ( .c(g6828), .b(g1377), .a(g5354) );
  and2_1361 AND2_193 ( .c(g8176), .b(g40), .a(n1173) );
  and2_1360 AND2_194 ( .c(g6830), .b(g1380), .a(g5354) );
  and2_1359 AND2_195 ( .c(g8005), .b(g7510), .a(n1253) );
  and2_1358 AND2_196 ( .c(g4099), .b(g770), .a(g3281) );
  and2_1357 AND2_197 ( .c(g11601), .b(g1351), .a(n1192) );
  and2_1356 AND2_198 ( .c(g11187), .b(g4727), .a(n1353) );
  and2_1355 AND2_199 ( .c(g6746), .b(g6228), .a(g5557) );
  and2_1354 AND2_200 ( .c(g6221), .b(g782), .a(g5598) );
  and2_1353 AND2_201 ( .c(g8765), .b(g8630), .a(g5151) );
  and2_1352 AND2_202 ( .c(g9622), .b(g1200), .a(g9111) );
  and2_1351 AND2_203 ( .c(g11143), .b(g10923), .a(n1164) );
  and2_1350 AND2_204 ( .c(g9904), .b(g9886), .a(g9676) );
  and2_1349 AND2_205 ( .c(g8733), .b(g8241), .a(n1384) );
  and3_41 AND3_8 ( .d(g8974), .c(n1260), .b(n1307), .a(n1281) );
  and2_1348 AND2_206 ( .c(g6624), .b(g348), .a(n1176) );
  and2_1347 AND2_207 ( .c(g11169), .b(g530), .a(n1346) );
  and2_1346 AND2_208 ( .c(g8073), .b(g709), .a(n1251) );
  and2_1345 AND2_209 ( .c(g9841), .b(g9706), .a(g9512) );
  and2_1344 AND2_210 ( .c(g5882), .b(g5592), .a(g3829) );
  and2_1343 AND2_211 ( .c(g8796), .b(g8645), .a(n1213) );
  and2_1342 AND2_212 ( .c(g11168), .b(g534), .a(n1346) );
  and2_1341 AND2_213 ( .c(g4269), .b(g1015), .a(n1371) );
  and2_1340 AND2_214 ( .c(g5271), .b(g727), .a(g3041) );
  and2_1339 AND2_215 ( .c(g10348), .b(n1219), .a(g109) );
  and2_1338 AND2_216 ( .c(g5611), .b(g1047), .a(n1371) );
  and2_1337 AND2_217 ( .c(g8069), .b(g673), .a(n1251) );
  and2_1336 AND2_218 ( .c(g9695), .b(g1567), .a(n1190) );
  and2_1335 AND2_219 ( .c(g10304), .b(g10001), .a(g8574) );
  and2_1334 AND2_220 ( .c(g8469), .b(g8305), .a(g7246) );
  and2_1333 AND2_221 ( .c(g4712), .b(g1071), .a(n1367) );
  and2_1332 AND2_222 ( .c(g6576), .b(g5762), .a(g3209) );
  and2_1331 AND2_223 ( .c(g10622), .b(g10496), .a(n1159) );
  and2_1330 AND2_224 ( .c(g11015), .b(g5217), .a(n1346) );
  and2_1329 AND2_225 ( .c(g5674), .b(g148), .a(g5361) );
  and2_1328 AND2_226 ( .c(g9359), .b(g1308), .a(n1328) );
  and2_1327 AND2_227 ( .c(g9223), .b(g48), .a(g8960) );
  and2_1326 AND2_228 ( .c(g11556), .b(g1786), .a(g11519) );
  and2_1325 AND2_229 ( .c(g9858), .b(g1595), .a(g9331) );
  and2_1324 AND2_230 ( .c(g5541), .b(g575), .a(n1391) );
  and2_1323 AND2_231 ( .c(g4534), .b(g363), .a(g3586) );
  and2_1322 AND2_232 ( .c(g6198), .b(g1499), .a(g5128) );
  and2_1321 AND2_233 ( .c(g6747), .b(n1151), .a(g5897) );
  and2_1320 AND2_234 ( .c(g6699), .b(g6177), .a(n1367) );
  and2_1319 AND2_235 ( .c(g6855), .b(n1145), .a(g6392) );
  and2_1318 AND2_236 ( .c(g3804), .b(g3098), .a(n1148) );
  and2_1317 AND2_237 ( .c(g5680), .b(g153), .a(g5361) );
  and2_1316 AND2_238 ( .c(g9642), .b(g981), .a(n1330) );
  and2_1315 AND2_239 ( .c(g5744), .b(g1528), .a(n1229) );
  and2_1314 AND2_240 ( .c(g10333), .b(n1219), .a(g109) );
  and2_1313 AND2_241 ( .c(g8399), .b(g5266), .a(g7101) );
  and2_1312 AND2_242 ( .c(g9447), .b(g1762), .a(n1329) );
  and2_1311 AND2_243 ( .c(g4903), .b(g1849), .a(n1288) );
  and2_1310 AND2_244 ( .c(g11178), .b(g516), .a(n1346) );
  and2_1309 AND2_245 ( .c(g8510), .b(g8414), .a(g7638) );
  and2_1308 AND2_246 ( .c(g8245), .b(g7062), .a(n1277) );
  and2_1307 AND2_247 ( .c(g6319), .b(g1296), .a(n1322) );
  and2_1306 AND2_248 ( .c(g11186), .b(g4722), .a(n1357) );
  and2_1305 AND2_249 ( .c(g3908), .b(g186), .a(n1386) );
  and2_1304 AND2_250 ( .c(g2951), .b(n1337), .a(g1681) );
  and2_1303 AND2_251 ( .c(g6352), .b(g278), .a(n1221) );
  and2_1302 AND2_252 ( .c(g9595), .b(g901), .a(g9205) );
  and2_1301 AND2_253 ( .c(g4831), .b(g810), .a(g4109) );
  and2_1300 AND2_254 ( .c(g5492), .b(g1654), .a(n1161) );
  and2_1299 AND2_255 ( .c(g9272), .b(g8934), .a(n1386) );
  and2_1298 AND2_256 ( .c(g10312), .b(g10019), .a(g8574) );
  and2_1297 AND2_257 ( .c(g6186), .b(g546), .a(n1372) );
  and2_1296 AND2_258 ( .c(g9612), .b(g971), .a(n1330) );
  and2_1295 AND2_259 ( .c(g9417), .b(g1738), .a(g9052) );
  and2_1294 AND2_260 ( .c(g9935), .b(g9914), .a(g9624) );
  and2_1293 AND2_261 ( .c(g8701), .b(n1234), .a(g8488) );
  and2_1292 AND2_262 ( .c(g10745), .b(g10658), .a(g3586) );
  and2_1291 AND2_263 ( .c(g11216), .b(g956), .a(n1177) );
  and2_1290 AND2_264 ( .c(g9328), .b(g8971), .a(g48) );
  and2_1289 AND2_265 ( .c(g11587), .b(g1327), .a(n1198) );
  and2_1288 AND2_266 ( .c(g6821), .b(g237), .a(g5354) );
  and2_1287 AND2_267 ( .c(g6325), .b(g1245), .a(n1322) );
  and2_1286 AND2_268 ( .c(g4560), .b(g431), .a(g109) );
  and2_1285 AND2_269 ( .c(g7368), .b(g5842), .a(g3880) );
  and2_1284 AND2_270 ( .c(g6083), .b(g552), .a(n1372) );
  and2_1283 AND2_271 ( .c(g6544), .b(g1227), .a(n1180) );
  and2_1282 AND2_272 ( .c(g5476), .b(g1615), .a(n1372) );
  and2_1281 AND2_273 ( .c(g7743), .b(g5838), .a(g3880) );
  and2_1280 AND2_274 ( .c(g4869), .b(g1083), .a(n1367) );
  and2_1279 AND2_275 ( .c(g5722), .b(g1598), .a(n1215) );
  and2_1278 AND2_276 ( .c(g6790), .b(g5813), .a(n1367) );
  and2_1277 AND2_277 ( .c(g8408), .b(g704), .a(n1211) );
  and2_1276 AND2_278 ( .c(g10761), .b(g10559), .a(g10558) );
  and2_1275 AND2_279 ( .c(g7734), .b(g5810), .a(g3880) );
  and2_1274 AND2_280 ( .c(g8136), .b(g7926), .a(n1253) );
  and2_1273 AND2_281 ( .c(g6187), .b(g5569), .a(n1111) );
  and2_1272 AND2_282 ( .c(g4752), .b(g401), .a(g109) );
  and2_1271 AND2_283 ( .c(g9902), .b(g9720), .a(n1321) );
  and2_1270 AND2_284 ( .c(g8768), .b(g8623), .a(g5151) );
  and2_1269 AND2_285 ( .c(g5500), .b(g1657), .a(n1161) );
  and2_1268 AND2_286 ( .c(g2496), .b(g374), .a(g369) );
  and2_1267 AND2_287 ( .c(g6756), .b(g3010), .a(g5877) );
  and3_40 AND3_9 ( .d(g8972), .c(n1271), .b(n1307), .a(n1281) );
  and2_1266 AND2_288 ( .c(g6622), .b(g336), .a(n1176) );
  and2_1265 AND2_289 ( .c(g11639), .b(g11612), .a(n1238) );
  and2_1264 AND2_290 ( .c(g9366), .b(g1311), .a(n1328) );
  and2_1263 AND2_291 ( .c(g11230), .b(n1334), .a(n1191) );
  and2_1262 AND2_292 ( .c(g10328), .b(n1220), .a(g109) );
  and2_1261 AND2_293 ( .c(g5024), .b(g1284), .a(g109) );
  and2_1260 AND2_294 ( .c(g4364), .b(g1215), .a(n1372) );
  and2_1259 AND2_295 ( .c(g9649), .b(g916), .a(g9205) );
  and2_1258 AND2_296 ( .c(g5795), .b(g1543), .a(n1229) );
  and2_1257 AND2_297 ( .c(g5737), .b(g1524), .a(n1229) );
  and2_1256 AND2_298 ( .c(g6841), .b(g1400), .a(g5354) );
  and2_1255 AND2_299 ( .c(g4054), .b(g1753), .a(n1206) );
  and2_1254 AND2_300 ( .c(g6345), .b(g5823), .a(n1366) );
  and2_1253 AND2_301 ( .c(g11391), .b(g11275), .a(n1237) );
  and2_1252 AND2_302 ( .c(g9851), .b(g296), .a(g9313) );
  and2_1251 AND2_303 ( .c(g6763), .b(g5802), .a(n1366) );
  and2_1250 AND2_304 ( .c(g4770), .b(g416), .a(g109) );
  and3_39 AND3_10 ( .d(I16142), .c(g10511), .b(g10509), .a(g10507) );
  and2_1249 AND2_305 ( .c(g9698), .b(g1571), .a(n1190) );
  and2_1248 AND2_306 ( .c(g4725), .b(g1032), .a(n1373) );
  and2_1247 AND2_307 ( .c(g5477), .b(g1887), .a(g3209) );
  and2_1246 AND2_308 ( .c(g9964), .b(g9954), .a(n1319) );
  and2_1245 AND2_309 ( .c(g5523), .b(g1663), .a(n1161) );
  and2_1244 AND2_310 ( .c(g4553), .b(g435), .a(g109) );
  and2_1243 AND2_311 ( .c(g8550), .b(g8402), .a(g7638) );
  and2_1242 AND2_312 ( .c(g8845), .b(g8611), .a(n1233) );
  and2_1241 AND2_313 ( .c(g2081), .b(g932), .a(g928) );
  and2_1240 AND2_314 ( .c(g6359), .b(g281), .a(n1221) );
  and2_1239 AND2_315 ( .c(g11586), .b(g1324), .a(n1198) );
  and2_1238 AND2_316 ( .c(g11007), .b(g5147), .a(n1346) );
  and2_1237 AND2_317 ( .c(g5104), .b(g1796), .a(n1202) );
  and2_1236 AND2_318 ( .c(g5099), .b(g4821), .a(g3829) );
  and2_1235 AND2_319 ( .c(g6757), .b(g143), .a(g5919) );
  and2_1234 AND2_320 ( .c(g5499), .b(g1627), .a(n1373) );
  and2_1233 AND2_321 ( .c(g4389), .b(g3529), .a(n1062) );
  and2_1232 AND2_322 ( .c(g6416), .b(g3497), .a(g5013) );
  and2_1231 AND2_323 ( .c(g9720), .b(g1546), .a(n1207) );
  and2_1230 AND2_324 ( .c(g4990), .b(g1444), .a(g4682) );
  and2_1229 AND2_325 ( .c(g9619), .b(g940), .a(n1326) );
  and4_15 AND4_1 ( .e(I6630), .d(n1333), .c(g1771), .b(g1776), .a(g1786) );
  and2_1228 AND2_326 ( .c(g6047), .b(n1129), .a(g4977) );
  and2_1227 AND2_327 ( .c(g9652), .b(g953), .a(n1324) );
  and3_38 AND3_11 ( .d(g10515), .c(g10505), .b(g10469), .a(I16142) );
  and2_1226 AND2_328 ( .c(g9843), .b(g9711), .a(g9519) );
  and2_1225 AND2_329 ( .c(g5273), .b(g1074), .a(n1161) );
  and2_1224 AND2_330 ( .c(g11465), .b(g11232), .a(g4421) );
  and2_1223 AND2_331 ( .c(g5044), .b(g4348), .a(g1918) );
  and2_1222 AND2_332 ( .c(g11237), .b(g4548), .a(n1355) );
  and2_1221 AND2_333 ( .c(g9834), .b(g9731), .a(g9785) );
  and2_1220 AND2_334 ( .c(g6654), .b(g363), .a(n1176) );
  and2_1219 AND2_335 ( .c(g5444), .b(g1041), .a(n1373) );
  and2_1218 AND2_336 ( .c(g3714), .b(n1337), .a(n1064) );
  and2_1217 AND2_337 ( .c(g11340), .b(g11285), .a(n1223) );
  and2_1216 AND2_338 ( .c(g9598), .b(g119), .a(n1323) );
  and2_1215 AND2_339 ( .c(g8097), .b(g5477), .a(g6740) );
  and2_1214 AND2_340 ( .c(g8726), .b(g8221), .a(n1384) );
  and2_1213 AND2_341 ( .c(g6880), .b(g4816), .a(n1267) );
  and2_1212 AND2_342 ( .c(g4338), .b(g1157), .a(g109) );
  and2_1211 AND2_343 ( .c(g5543), .b(g2979), .a(n1277) );
  and3_37 AND3_12 ( .d(g8960), .c(n1271), .b(n1307), .a(n1266) );
  and2_1210 AND2_344 ( .c(g4109), .b(g806), .a(g3287) );
  and2_1209 AND2_345 ( .c(g10759), .b(g10557), .a(g10556) );
  and2_1208 AND2_346 ( .c(g9938), .b(g9917), .a(n1320) );
  and2_1207 AND2_347 ( .c(g10758), .b(g10652), .a(n1366) );
  and2_1206 AND2_348 ( .c(g4759), .b(g406), .a(g109) );
  and2_1205 AND2_349 ( .c(g9909), .b(g9891), .a(n1327) );
  and2_1204 AND2_350 ( .c(g7127), .b(g6663), .a(n1106) );
  and2_1203 AND2_351 ( .c(g11165), .b(g476), .a(n1346) );
  and2_1202 AND2_352 ( .c(g6234), .b(g1424), .a(g5151) );
  and2_1201 AND2_353 ( .c(g6328), .b(g1260), .a(n1322) );
  and2_1200 AND2_354 ( .c(g8401), .b(g677), .a(n1211) );
  and2_1199 AND2_355 ( .c(g11006), .b(g5125), .a(n1346) );
  and2_1198 AND2_356 ( .c(g4865), .b(g1080), .a(n1366) );
  and2_1197 AND2_357 ( .c(g4715), .b(g1077), .a(n1366) );
  and3_36 AND3_13 ( .d(g4604), .c(g3056), .b(g3753), .a(g2325) );
  and2_1196 AND2_358 ( .c(g5513), .b(g1675), .a(n1373) );
  and2_1195 AND2_359 ( .c(g11222), .b(g965), .a(n1177) );
  and2_1194 AND2_360 ( .c(g4498), .b(g1145), .a(g109) );
  and2_1193 AND2_361 ( .c(g6554), .b(g96), .a(n1316) );
  and2_1192 AND2_362 ( .c(g7732), .b(g5803), .a(g3880) );
  and2_1191 AND2_363 ( .c(g9586), .b(g1346), .a(n1328) );
  and3_35 AND3_14 ( .d(g5178), .c(n1084), .b(g4401), .a(g4104) );
  and2_1190 AND2_364 ( .c(g4584), .b(n1282), .a(g1857) );
  and2_1189 AND2_365 ( .c(g7472), .b(n1384), .a(g61) );
  and2_1188 AND2_366 ( .c(g11253), .b(g981), .a(n1169) );
  and2_1187 AND2_367 ( .c(g5182), .b(g1240), .a(g109) );
  and2_1186 AND2_368 ( .c(g9860), .b(g1598), .a(g9331) );
  and2_1185 AND2_369 ( .c(g8703), .b(n1234), .a(g8488) );
  and2_1184 AND2_370 ( .c(g11600), .b(g1346), .a(n1192) );
  and2_1183 AND2_371 ( .c(g9710), .b(g1586), .a(n1190) );
  and2_1182 AND2_372 ( .c(g9645), .b(g1203), .a(g9111) );
  and2_1181 AND2_373 ( .c(g11236), .b(g4537), .a(n1353) );
  and2_1180 AND2_374 ( .c(g4162), .b(g3106), .a(g1845) );
  and2_1179 AND2_375 ( .c(g6090), .b(g553), .a(n1374) );
  and2_1178 AND2_376 ( .c(g9691), .b(g269), .a(n1171) );
  and2_1177 AND2_377 ( .c(g11372), .b(g11316), .a(n1223) );
  and2_1176 AND2_378 ( .c(g6823), .b(g1368), .a(g5354) );
  and2_1175 AND2_379 ( .c(g11175), .b(g501), .a(n1346) );
  and2_1174 AND2_380 ( .c(g8068), .b(g664), .a(n1251) );
  and2_1173 AND2_381 ( .c(g9607), .b(g12), .a(n1323) );
  and2_1172 AND2_382 ( .c(g9962), .b(g9952), .a(n1319) );
  and2_1171 AND2_383 ( .c(g6348), .b(g296), .a(n1221) );
  and2_1170 AND2_384 ( .c(g9659), .b(g956), .a(n1324) );
  and2_1169 AND2_385 ( .c(g9358), .b(g1318), .a(n1325) );
  and2_1168 AND2_386 ( .c(g3104), .b(I6316), .a(I6317) );
  and2_1167 AND2_387 ( .c(g4486), .b(g1711), .a(n1374) );
  and2_1166 AND2_388 ( .c(g9587), .b(g892), .a(g8995) );
  and2_1165 AND2_389 ( .c(g5632), .b(g1636), .a(n1390) );
  and2_1164 AND2_390 ( .c(g9111), .b(g8965), .a(g48) );
  and2_1163 AND2_391 ( .c(g4881), .b(g991), .a(n1374) );
  and2_1162 AND2_392 ( .c(g11209), .b(g10712), .a(n1224) );
  and2_1161 AND2_393 ( .c(g8848), .b(g8715), .a(n1233) );
  and2_1160 AND2_394 ( .c(g4070), .b(g3263), .a(n1125) );
  and2_1159 AND2_395 ( .c(g6463), .b(g48), .a(n1306) );
  and2_1158 AND2_396 ( .c(g8699), .b(n1234), .a(g8488) );
  and4_14 AND4_2 ( .e(I5689), .d(g1419), .c(g1424), .b(g1428), .a(g1432) );
  and2_1157 AND2_397 ( .c(g7820), .b(g1896), .a(n1257) );
  and2_1156 AND2_398 ( .c(g11021), .b(g448), .a(n1347) );
  and2_1155 AND2_399 ( .c(g5917), .b(g1044), .a(g85) );
  and2_1154 AND2_400 ( .c(g6619), .b(g49), .a(n1176) );
  and2_1153 AND2_401 ( .c(g6318), .b(g1300), .a(n1322) );
  and2_1152 AND2_402 ( .c(g6872), .b(g1896), .a(g6003) );
  and2_1151 AND2_403 ( .c(g11320), .b(g11201), .a(n1208) );
  and2_1150 AND2_404 ( .c(g10514), .b(g10489), .a(n1159) );
  and2_1149 AND2_405 ( .c(g4006), .b(g201), .a(n1386) );
  and2_1148 AND2_406 ( .c(g9853), .b(g299), .a(g9313) );
  and2_1147 AND2_407 ( .c(g11274), .b(g4771), .a(n1344) );
  and2_1146 AND2_408 ( .c(g6193), .b(g1419), .a(g5151) );
  and2_1145 AND2_409 ( .c(g8119), .b(g5526), .a(g6740) );
  and2_1144 AND2_410 ( .c(g9420), .b(g1747), .a(n1329) );
  and2_1143 AND2_411 ( .c(g5233), .b(g1791), .a(g4492) );
  and2_1142 AND2_412 ( .c(g7581), .b(g7092), .a(n1240) );
  and2_1141 AND2_413 ( .c(g6549), .b(g95), .a(n1316) );
  and2_1140 AND2_414 ( .c(g11464), .b(g11231), .a(g4421) );
  and2_1139 AND2_415 ( .c(g4801), .b(g516), .a(g109) );
  and2_1138 AND2_416 ( .c(g6834), .b(g1365), .a(g5354) );
  and2_1137 AND2_417 ( .c(g4487), .b(g1718), .a(n1374) );
  and2_1136 AND2_418 ( .c(g2939), .b(n1337), .a(g1687) );
  and2_1135 AND2_419 ( .c(g7060), .b(g6739), .a(g3041) );
  and2_1134 AND2_420 ( .c(g5770), .b(g3585), .a(g5128) );
  and2_1133 AND2_421 ( .c(g5725), .b(g1580), .a(n1215) );
  and2_1132 AND2_422 ( .c(g11641), .b(g11615), .a(n1238) );
  and2_1131 AND2_423 ( .c(g2544), .b(g1341), .a(g1336) );
  and2_1130 AND2_424 ( .c(g11292), .b(g11252), .a(n1208) );
  and2_1129 AND2_425 ( .c(g5532), .b(g1681), .a(n1375) );
  and2_1128 AND2_426 ( .c(g11153), .b(g3771), .a(g10788) );
  and2_1127 AND2_427 ( .c(g9905), .b(g9872), .a(g9680) );
  and2_1126 AND2_428 ( .c(g7739), .b(g5820), .a(g3880) );
  and2_1125 AND2_429 ( .c(g6321), .b(g1284), .a(n1322) );
  and2_1124 AND2_430 ( .c(g8386), .b(g5257), .a(g7101) );
  and3_34 AND3_15 ( .d(g8975), .c(n1268), .b(n1307), .a(n1281) );
  and2_1123 AND2_431 ( .c(g2306), .b(g1223), .a(g1218) );
  and2_1122 AND2_432 ( .c(g6625), .b(g1218), .a(n1180) );
  and2_1121 AND2_433 ( .c(g7937), .b(g5274), .a(n1366) );
  and2_1120 AND2_434 ( .c(g10788), .b(g8303), .a(n1347) );
  and2_1119 AND2_435 ( .c(g10325), .b(n1232), .a(g109) );
  and2_1118 AND2_436 ( .c(g8170), .b(g36), .a(n1173) );
  and2_1117 AND2_437 ( .c(g5706), .b(g1574), .a(n1215) );
  and2_1116 AND2_438 ( .c(g2756), .b(g936), .a(g2081) );
  and2_1115 AND2_439 ( .c(g8821), .b(g8643), .a(n1233) );
  and2_1114 AND2_440 ( .c(g10946), .b(g5225), .a(n1347) );
  and2_1113 AND2_441 ( .c(g4169), .b(g1806), .a(n1103) );
  and2_1112 AND2_442 ( .c(g5029), .b(g1077), .a(n1161) );
  and2_1111 AND2_443 ( .c(g11164), .b(g3513), .a(n1347) );
  and2_1110 AND2_444 ( .c(g4007), .b(g1771), .a(g2276) );
  and2_1109 AND2_445 ( .c(g4059), .b(g1756), .a(n1206) );
  and2_1108 AND2_446 ( .c(g4868), .b(g1027), .a(n1375) );
  and2_1107 AND2_447 ( .c(g5675), .b(g131), .a(g5361) );
  and2_1106 AND2_448 ( .c(g4718), .b(g650), .a(n1089) );
  and2_1105 AND2_449 ( .c(g10682), .b(g10381), .a(g3863) );
  and2_1104 AND2_450 ( .c(g6687), .b(g92), .a(n1316) );
  and2_1103 AND2_451 ( .c(g7704), .b(g682), .a(g6488) );
  and2_1102 AND2_452 ( .c(g4582), .b(g525), .a(g109) );
  and2_1101 AND2_453 ( .c(g4261), .b(g1019), .a(n1375) );
  and2_1100 AND2_454 ( .c(g3422), .b(g225), .a(n1386) );
  and2_1099 AND2_455 ( .c(g5745), .b(g1549), .a(n1229) );
  and2_1098 AND2_456 ( .c(g8387), .b(g5258), .a(g7101) );
  and2_1097 AND2_457 ( .c(g7954), .b(g49), .a(n1383) );
  and2_1096 AND2_458 ( .c(g11283), .b(g4804), .a(n1352) );
  and2_1095 AND2_459 ( .c(g8461), .b(g8298), .a(g7246) );
  and2_1094 AND2_460 ( .c(g10760), .b(g10555), .a(g10554) );
  and2_1093 AND2_461 ( .c(g11492), .b(g11480), .a(n1322) );
  and3_33 AND3_16 ( .d(g7032), .c(g109), .b(g6626), .a(n1295) );
  and2_1092 AND2_462 ( .c(g8756), .b(n1231), .a(g8451) );
  and2_1091 AND2_463 ( .c(g9151), .b(g8967), .a(g48) );
  and2_1090 AND2_464 ( .c(g6341), .b(g272), .a(n1221) );
  and2_1089 AND2_465 ( .c(g10506), .b(g10007), .a(n1337) );
  and2_1088 AND2_466 ( .c(g9648), .b(g16), .a(n1323) );
  and2_1087 AND2_467 ( .c(g7453), .b(n1384), .a(g52) );
  and2_1086 AND2_468 ( .c(g6525), .b(g5995), .a(n1083) );
  and2_1085 AND2_469 ( .c(g6645), .b(g67), .a(n1176) );
  and2_1084 AND2_470 ( .c(g5707), .b(g1595), .a(n1215) );
  and2_1083 AND2_471 ( .c(g8046), .b(g7548), .a(g5128) );
  and2_1082 AND2_472 ( .c(g11091), .b(g833), .a(g10950) );
  and2_1081 AND2_473 ( .c(g11174), .b(g496), .a(n1347) );
  and2_1080 AND2_474 ( .c(g9010), .b(g48), .a(g8930) );
  and2_1079 AND2_475 ( .c(g8403), .b(g5276), .a(g7101) );
  and2_1078 AND2_476 ( .c(g5201), .b(g1250), .a(g109) );
  and2_1077 AND2_477 ( .c(g8841), .b(g8605), .a(n1233) );
  and2_1076 AND2_478 ( .c(g6879), .b(g1914), .a(g6003) );
  and2_1075 AND2_479 ( .c(g8763), .b(n1231), .a(g8451) );
  and2_1074 AND2_480 ( .c(g4502), .b(n1103), .a(g1707) );
  and2_1073 AND2_481 ( .c(g9839), .b(g9702), .a(g9742) );
  and2_1072 AND2_482 ( .c(g6358), .b(g5841), .a(n1366) );
  and2_1071 AND2_483 ( .c(g5575), .b(g1618), .a(n1390) );
  and2_1070 AND2_484 ( .c(g4940), .b(n1070), .a(n1286) );
  and2_1069 AND2_485 ( .c(g8107), .b(g5502), .a(g6740) );
  and2_1068 AND2_486 ( .c(g10240), .b(g9974), .a(g8574) );
  and2_1067 AND2_487 ( .c(g11192), .b(g4759), .a(n1344) );
  and2_1066 AND2_488 ( .c(g9618), .b(g910), .a(g9205) );
  and2_1065 AND2_489 ( .c(g5539), .b(g1684), .a(n1375) );
  and2_1064 AND2_490 ( .c(g8416), .b(g731), .a(n1211) );
  and2_1063 AND2_491 ( .c(g9693), .b(g275), .a(n1171) );
  and2_1062 AND2_492 ( .c(g11553), .b(g1771), .a(g11519) );
  and2_1061 AND2_493 ( .c(g8047), .b(g7557), .a(g5919) );
  and2_1060 AND2_494 ( .c(g5268), .b(g1098), .a(n1161) );
  and2_1059 AND2_495 ( .c(g9555), .b(g9107), .a(n1386) );
  and2_1058 AND2_496 ( .c(g6180), .b(g1453), .a(g5128) );
  and2_1057 AND2_497 ( .c(g6832), .b(g1383), .a(g5354) );
  and2_1056 AND2_498 ( .c(g10633), .b(g10381), .a(g3829) );
  and2_1055 AND2_499 ( .c(g7894), .b(g5317), .a(n1390) );
  and2_1054 AND2_500 ( .c(g8654), .b(g8266), .a(n1366) );
  and2_1053 AND2_501 ( .c(g9621), .b(g1179), .a(g9125) );
  and2_1052 AND2_502 ( .c(g6794), .b(g5819), .a(n1366) );
  and2_1051 AND2_503 ( .c(g9313), .b(g8876), .a(g48) );
  and2_1050 AND2_504 ( .c(g4883), .b(g248), .a(n1386) );
  and2_1049 AND2_505 ( .c(g3412), .b(g219), .a(n1386) );
  and2_1048 AND2_506 ( .c(g7661), .b(g7127), .a(n1127) );
  and3_32 AND3_17 ( .d(g2800), .c(n1130), .b(n1099), .a(g591) );
  and2_1047 AND2_507 ( .c(g3389), .b(g207), .a(n1386) );
  and2_1046 AND2_508 ( .c(g3706), .b(n1334), .a(g3268) );
  and2_1045 AND2_509 ( .c(g9908), .b(n1182), .a(n1327) );
  and2_1044 AND2_510 ( .c(g3429), .b(g231), .a(n1386) );
  and2_1043 AND2_511 ( .c(g6628), .b(g351), .a(n1176) );
  and2_1042 AND2_512 ( .c(g5470), .b(g1044), .a(n1376) );
  and2_1041 AND2_513 ( .c(g7526), .b(n1384), .a(g73) );
  and2_1040 AND2_514 ( .c(g5897), .b(g2204), .a(g5354) );
  and2_1039 AND2_515 ( .c(g5025), .b(g1482), .a(g4640) );
  and2_1038 AND2_516 ( .c(g6204), .b(n1280), .a(g4921) );
  and2_1037 AND2_517 ( .c(g4048), .b(g1750), .a(n1206) );
  and3_31 AND3_18 ( .d(g8935), .c(n1250), .b(n1307), .a(n1274) );
  and2_1036 AND2_518 ( .c(g3281), .b(g766), .a(g2525) );
  and2_1035 AND2_519 ( .c(g9593), .b(g898), .a(g9205) );
  and2_1034 AND2_520 ( .c(g4827), .b(g213), .a(n1386) );
  and2_1033 AND2_521 ( .c(g10701), .b(g10501), .a(g10500) );
  and2_1032 AND2_522 ( .c(g10777), .b(g10733), .a(n1366) );
  and2_1031 AND2_523 ( .c(g8130), .b(g1936), .a(n1210) );
  and2_1030 AND2_524 ( .c(g9965), .b(g9955), .a(n1319) );
  and2_1029 AND2_525 ( .c(g3684), .b(g1710), .a(n1366) );
  and2_1028 AND2_526 ( .c(g11213), .b(g947), .a(n1177) );
  and2_1027 AND2_527 ( .c(g5006), .b(g1462), .a(g4640) );
  and2_1026 AND2_528 ( .c(g9933), .b(g9912), .a(g9624) );
  and2_1025 AND2_529 ( .c(g8554), .b(g8407), .a(g7638) );
  and2_1024 AND2_530 ( .c(g9641), .b(g913), .a(g9205) );
  and2_1023 AND2_531 ( .c(g6123), .b(g3662), .a(n1286) );
  and2_1022 AND2_532 ( .c(g6323), .b(g1235), .a(n1322) );
  and2_1021 AND2_533 ( .c(g10766), .b(g10646), .a(n1366) );
  and2_1020 AND2_534 ( .c(g6666), .b(g89), .a(n1316) );
  and2_1019 AND2_535 ( .c(g4994), .b(g1504), .a(g4640) );
  and2_1018 AND2_536 ( .c(g5755), .b(g5103), .a(g5354) );
  and2_1017 AND2_537 ( .c(g11592), .b(g3717), .a(g11561) );
  and2_1016 AND2_538 ( .c(g6351), .b(n1306), .a(g48) );
  and2_1015 AND2_539 ( .c(g6875), .b(g1905), .a(g6003) );
  and2_1014 AND2_540 ( .c(g4816), .b(g4070), .a(n1120) );
  and2_1013 AND2_541 ( .c(g9658), .b(g947), .a(n1330) );
  and2_1012 AND2_542 ( .c(g6530), .b(g6207), .a(g3829) );
  and2_1011 AND2_543 ( .c(g8366), .b(g8199), .a(g7265) );
  and2_1010 AND2_544 ( .c(g9835), .b(g9735), .a(g9785) );
  and2_1009 AND2_545 ( .c(g6655), .b(g88), .a(n1316) );
  and3_30 AND3_19 ( .d(g5445), .c(n1295), .b(g3875), .a(g109) );
  and2_1008 AND2_546 ( .c(g5173), .b(n1338), .a(n1235) );
  and2_1007 AND2_547 ( .c(g7970), .b(g7384), .a(n1245) );
  and2_1006 AND2_548 ( .c(g3098), .b(n1137), .a(n1135) );
  and2_1005 AND2_549 ( .c(g5491), .b(g1624), .a(n1376) );
  and2_1004 AND2_550 ( .c(g9271), .b(n1385), .a(g8949) );
  and2_1003 AND2_551 ( .c(g11152), .b(g369), .a(n1163) );
  and2_1002 AND2_552 ( .c(g9611), .b(g936), .a(n1326) );
  and2_1001 AND2_553 ( .c(g6410), .b(g2804), .a(g5013) );
  and2_1000 AND2_554 ( .c(g10451), .b(n1170), .a(n1071) );
  and2_999 AND2_555 ( .c(g4397), .b(n1244), .a(g639) );
  and2_998 AND2_556 ( .c(g7224), .b(g5398), .a(n1276) );
  and2_997 AND2_557 ( .c(g5602), .b(g1624), .a(n1390) );
  and2_996 AND2_558 ( .c(g4421), .b(n1144), .a(g750) );
  and2_995 AND2_559 ( .c(g6884), .b(g5569), .a(n1267) );
  and2_994 AND2_560 ( .c(g6839), .b(g1397), .a(g5354) );
  and2_993 AND2_561 ( .c(g8698), .b(n1234), .a(g8488) );
  and3_29 AND3_20 ( .d(g8964), .c(n1259), .b(n1307), .a(n1274) );
  and2_992 AND2_562 ( .c(g8260), .b(g940), .a(n1209) );
  and2_991 AND2_563 ( .c(g11413), .b(g11217), .a(g10522) );
  and2_990 AND2_564 ( .c(g4950), .b(g1415), .a(g4682) );
  and2_989 AND2_565 ( .c(g5535), .b(g572), .a(n1390) );
  and2_988 AND2_566 ( .c(g7277), .b(g6772), .a(g731) );
  and2_987 AND2_567 ( .c(g8463), .b(g8301), .a(g7246) );
  and2_986 AND2_568 ( .c(g3268), .b(n1335), .a(g2511) );
  and2_985 AND2_569 ( .c(g10785), .b(g10728), .a(n1202) );
  and2_984 AND2_570 ( .c(g6618), .b(g658), .a(g5557) );
  and2_983 AND2_571 ( .c(g6235), .b(g569), .a(n1376) );
  and2_982 AND2_572 ( .c(g10950), .b(g10788), .a(g6355) );
  and2_981 AND2_573 ( .c(g4723), .b(g3626), .a(g627) );
  and2_980 AND2_574 ( .c(g8720), .b(g8206), .a(n1384) );
  and2_979 AND2_575 ( .c(g6693), .b(g93), .a(n1316) );
  and2_978 AND2_576 ( .c(g11020), .b(g452), .a(n1347) );
  and2_977 AND2_577 ( .c(g11583), .b(g1314), .a(n1198) );
  and2_976 AND2_578 ( .c(g8118), .b(g1900), .a(n1210) );
  and2_975 AND2_579 ( .c(g8167), .b(g33), .a(n1173) );
  and2_974 AND2_580 ( .c(g6334), .b(g1389), .a(g5354) );
  and2_973 AND2_581 ( .c(g7892), .b(g5308), .a(n1391) );
  and2_972 AND2_582 ( .c(g8652), .b(g8264), .a(n1365) );
  and2_971 AND2_583 ( .c(g5721), .b(g1577), .a(n1215) );
  and2_970 AND2_584 ( .c(g10367), .b(g10362), .a(n1071) );
  and2_969 AND2_585 ( .c(g9901), .b(g9719), .a(n1321) );
  and2_968 AND2_586 ( .c(g6792), .b(g290), .a(n1221) );
  and2_967 AND2_587 ( .c(g11282), .b(g4801), .a(n1354) );
  and2_966 AND2_588 ( .c(g7945), .b(g67), .a(n1383) );
  and3_28 AND3_21 ( .d(g8971), .c(n1284), .b(n1307), .a(n1281) );
  and2_965 AND2_589 ( .c(g11302), .b(g4582), .a(n1353) );
  and2_964 AND2_590 ( .c(g4585), .b(g521), .a(g109) );
  and2_963 AND2_591 ( .c(g6621), .b(g52), .a(n1176) );
  and2_962 AND2_592 ( .c(g5502), .b(g1932), .a(g3209) );
  and2_961 AND2_593 ( .c(g11105), .b(g3634), .a(g10937) );
  and2_960 AND2_594 ( .c(g7709), .b(g5942), .a(n1277) );
  and2_959 AND2_595 ( .c(g8598), .b(g8471), .a(g7246) );
  and2_958 AND2_596 ( .c(g7140), .b(g5221), .a(n1199) );
  and2_957 AND2_597 ( .c(g9600), .b(g904), .a(g9205) );
  and2_956 AND2_598 ( .c(g9864), .b(g1604), .a(g9331) );
  and2_955 AND2_599 ( .c(g11640), .b(g11613), .a(n1238) );
  and2_954 AND2_600 ( .c(g5188), .b(g798), .a(g794) );
  and2_953 AND2_601 ( .c(g7435), .b(g7260), .a(n1267) );
  and2_952 AND2_602 ( .c(g7876), .b(g5278), .a(n1391) );
  and2_951 AND2_603 ( .c(g5030), .b(g1280), .a(g109) );
  and2_950 AND2_604 ( .c(g4058), .b(g1791), .a(g2276) );
  and2_949 AND2_605 ( .c(g6776), .b(g5809), .a(n1365) );
  and2_948 AND2_606 ( .c(g4890), .b(g630), .a(n1263) );
  and2_947 AND2_607 ( .c(g2525), .b(g762), .a(g758) );
  and2_946 AND2_608 ( .c(g10301), .b(n1224), .a(g10025) );
  and2_945 AND2_609 ( .c(g4505), .b(g354), .a(g3586) );
  and2_944 AND2_610 ( .c(g9623), .b(g17), .a(n1323) );
  and2_943 AND2_611 ( .c(g10739), .b(n1294), .a(n1298) );
  and2_942 AND2_612 ( .c(g11027), .b(g391), .a(n1347) );
  and2_941 AND2_613 ( .c(g10738), .b(g10599), .a(n1365) );
  and2_940 AND2_614 ( .c(g8687), .b(g8558), .a(g7638) );
  and2_939 AND2_615 ( .c(g6360), .b(g302), .a(n1221) );
  and2_938 AND2_616 ( .c(g9871), .b(g1564), .a(g9324) );
  and2_937 AND2_617 ( .c(g5108), .b(g1801), .a(n1202) );
  and2_936 AND2_618 ( .c(g11248), .b(g976), .a(n1169) );
  and2_935 AND2_619 ( .c(g4992), .b(g1407), .a(g4682) );
  and2_934 AND2_620 ( .c(g11552), .b(n1333), .a(g11519) );
  and2_933 AND2_621 ( .c(g9651), .b(g944), .a(n1330) );
  and2_932 AND2_622 ( .c(g11204), .b(g971), .a(n1169) );
  and2_931 AND2_623 ( .c(g7824), .b(g1932), .a(n1257) );
  and2_930 AND2_624 ( .c(g4480), .b(g1133), .a(g109) );
  and2_929 AND2_625 ( .c(g6179), .b(g5115), .a(g5354) );
  and2_928 AND2_626 ( .c(g8710), .b(n1234), .a(g8488) );
  and2_927 AND2_627 ( .c(g7590), .b(g7102), .a(n1240) );
  and2_926 AND2_628 ( .c(g9384), .b(g968), .a(n1324) );
  and2_925 AND2_629 ( .c(g3407), .b(g2561), .a(g109) );
  and2_924 AND2_630 ( .c(g9838), .b(g9700), .a(g9754) );
  and2_923 AND2_631 ( .c(g3718), .b(g192), .a(n1386) );
  and2_922 AND2_632 ( .c(g10661), .b(g10594), .a(n1365) );
  and2_921 AND2_633 ( .c(g11380), .b(g11321), .a(n1223) );
  and3_27 AND3_22 ( .d(g8879), .c(n1283), .b(n1307), .a(n1281) );
  and2_920 AND2_634 ( .c(g7930), .b(g7621), .a(n1083) );
  and3_26 AND3_23 ( .d(g8962), .c(n1268), .b(n1307), .a(n1266) );
  and2_919 AND2_635 ( .c(g10715), .b(g2272), .a(n1299) );
  and2_918 AND2_636 ( .c(g8659), .b(g8269), .a(n1365) );
  and2_917 AND2_637 ( .c(g3015), .b(n1132), .a(n1301) );
  and2_916 AND2_638 ( .c(g9643), .b(g950), .a(n1324) );
  and2_915 AND2_639 ( .c(g9205), .b(g48), .a(g8957) );
  and2_914 AND2_640 ( .c(g5538), .b(g1669), .a(n1161) );
  and2_913 AND2_641 ( .c(g4000), .b(g1744), .a(n1206) );
  and2_912 AND2_642 ( .c(g4126), .b(g1786), .a(n1103) );
  and2_911 AND2_643 ( .c(g4400), .b(g4088), .a(g3829) );
  and2_910 AND2_644 ( .c(g2794), .b(I5886), .a(I5887) );
  and2_909 AND2_645 ( .c(g4760), .b(g486), .a(g109) );
  and2_908 AND2_646 ( .c(g6238), .b(g572), .a(n1376) );
  and2_907 AND2_647 ( .c(g10784), .b(g10727), .a(n1202) );
  and2_906 AND2_648 ( .c(g8174), .b(g38), .a(n1173) );
  and2_905 AND2_649 ( .c(g6332), .b(g1374), .a(g5354) );
  and2_904 AND2_650 ( .c(g5067), .b(g305), .a(n1196) );
  and2_903 AND2_651 ( .c(g5418), .b(g1512), .a(n1389) );
  and2_902 AND2_652 ( .c(g10297), .b(n1224), .a(g10001) );
  and2_901 AND2_653 ( .c(g6353), .b(g299), .a(n1221) );
  and2_900 AND2_654 ( .c(g11026), .b(g386), .a(n1347) );
  and2_899 AND2_655 ( .c(g11212), .b(g944), .a(n1177) );
  and2_898 AND2_656 ( .c(g6744), .b(g4828), .a(g5557) );
  and2_897 AND2_657 ( .c(g5493), .b(g1923), .a(g3209) );
  and2_896 AND2_658 ( .c(g10671), .b(g10411), .a(n1224) );
  and2_895 AND2_659 ( .c(g4383), .b(g2517), .a(g3829) );
  and2_894 AND2_660 ( .c(g5256), .b(g4297), .a(g627) );
  and2_893 AND2_661 ( .c(g4220), .b(g105), .a(n1377) );
  and2_892 AND2_662 ( .c(g8380), .b(g8252), .a(g3209) );
  and2_891 AND2_663 ( .c(g7071), .b(g5030), .a(n1199) );
  and2_890 AND2_664 ( .c(g4779), .b(g501), .a(g109) );
  and2_889 AND2_665 ( .c(g9613), .b(g1176), .a(g9125) );
  and2_888 AND2_666 ( .c(g7705), .b(g5935), .a(n1286) );
  and2_887 AND2_667 ( .c(g9269), .b(g8933), .a(n1386) );
  and2_886 AND2_668 ( .c(g5181), .b(g806), .a(g802) );
  and2_885 AND2_669 ( .c(g4977), .b(n1164), .a(n1322) );
  and2_884 AND2_670 ( .c(g7948), .b(g70), .a(n1383) );
  and2_883 AND2_671 ( .c(g11149), .b(g324), .a(n1353) );
  and2_882 AND2_672 ( .c(g9862), .b(g1601), .a(g9331) );
  and2_881 AND2_673 ( .c(g11387), .b(g11077), .a(n1389) );
  and2_880 AND2_674 ( .c(g7955), .b(g76), .a(n1383) );
  and2_879 AND2_675 ( .c(g4161), .b(g1801), .a(n1103) );
  and2_878 AND2_676 ( .c(g11148), .b(g2321), .a(g10788) );
  and2_877 AND2_677 ( .c(g9712), .b(g1528), .a(n1207) );
  and2_876 AND2_678 ( .c(g8931), .b(g8642), .a(g41) );
  and2_875 AND2_679 ( .c(g11097), .b(g378), .a(n1163) );
  and3_25 AND3_24 ( .d(g5421), .c(n1295), .b(g109), .a(g3819) );
  and2_874 AND2_680 ( .c(g11104), .b(g2963), .a(g10937) );
  and2_873 AND2_681 ( .c(g5263), .b(g709), .a(g3041) );
  and2_872 AND2_682 ( .c(g6092), .b(g1059), .a(g85) );
  and2_871 AND2_683 ( .c(g4999), .b(g1499), .a(g4640) );
  and4_13 AND4_3 ( .e(I6338), .d(n1105), .c(n1080), .b(n1063), .a(n1085) );
  and3_24 AND3_25 ( .d(g7409), .c(g4976), .b(g632), .a(g6858) );
  and2_870 AND2_684 ( .c(g4103), .b(g1771), .a(n1103) );
  and4_12 AND4_4 ( .e(I6309), .d(n1085), .c(n1063), .b(n1080), .a(n1105) );
  and2_869 AND2_685 ( .c(g6580), .b(g1801), .a(g5944) );
  and2_868 AND2_686 ( .c(g5631), .b(g1056), .a(n1377) );
  and2_867 AND2_687 ( .c(g9414), .b(g1730), .a(g9052) );
  and2_866 AND2_688 ( .c(g9660), .b(g1188), .a(g9125) );
  and2_865 AND2_689 ( .c(g9946), .b(g9926), .a(n1321) );
  and2_864 AND2_690 ( .c(g5257), .b(g691), .a(g3041) );
  and2_863 AND2_691 ( .c(g4732), .b(g391), .a(g109) );
  and2_862 AND2_692 ( .c(g3108), .b(I6330), .a(I6331) );
  and2_861 AND2_693 ( .c(g4753), .b(g481), .a(g109) );
  and2_860 AND2_694 ( .c(g9903), .b(g9885), .a(g9673) );
  and2_859 AND2_695 ( .c(g10625), .b(g10454), .a(n1159) );
  and2_858 AND2_696 ( .c(g5605), .b(g4828), .a(g704) );
  and2_857 AND2_697 ( .c(g6623), .b(g55), .a(n1176) );
  and2_856 AND2_698 ( .c(g11228), .b(n1335), .a(n1191) );
  and2_855 AND2_699 ( .c(g11011), .b(n1051), .a(g10809) );
  and2_854 AND2_700 ( .c(g6889), .b(g1941), .a(g6003) );
  and2_853 AND2_701 ( .c(g8040), .b(g7523), .a(g5128) );
  and2_852 AND2_702 ( .c(g7822), .b(g1914), .a(n1257) );
  and2_851 AND2_703 ( .c(g8123), .b(g1918), .a(n1210) );
  and2_850 AND2_704 ( .c(g11582), .b(g1311), .a(n1198) );
  and2_849 AND2_705 ( .c(g4316), .b(n1134), .a(g3400) );
  and2_848 AND2_706 ( .c(g10969), .b(g3625), .a(g10809) );
  and2_847 AND2_707 ( .c(g5041), .b(n1278), .a(g4401) );
  and2_846 AND2_708 ( .c(g9335), .b(g8975), .a(g48) );
  and2_845 AND2_709 ( .c(g9831), .b(g9727), .a(g9785) );
  and2_844 AND2_710 ( .c(g4565), .b(g534), .a(g109) );
  and2_843 AND2_711 ( .c(g9422), .b(g1750), .a(n1329) );
  and2_842 AND2_712 ( .c(g8648), .b(g4588), .a(g8511) );
  and3_23 AND3_26 ( .d(g8875), .c(n1259), .b(n1307), .a(n1281) );
  and2_841 AND2_713 ( .c(g5168), .b(g1512), .a(n1377) );
  and2_840 AND2_714 ( .c(g7895), .b(g7503), .a(n1253) );
  and2_839 AND2_715 ( .c(g8655), .b(g8267), .a(n1365) );
  and2_838 AND2_716 ( .c(g3396), .b(g213), .a(n1386) );
  and2_837 AND2_717 ( .c(g4914), .b(g1062), .a(n1377) );
  and2_836 AND2_718 ( .c(g9947), .b(g9927), .a(n1321) );
  and2_835 AND2_719 ( .c(g5772), .b(g1555), .a(n1229) );
  and2_834 AND2_720 ( .c(g6838), .b(g192), .a(g5354) );
  and2_833 AND2_721 ( .c(g5531), .b(g1666), .a(n1161) );
  and2_832 AND2_722 ( .c(g6795), .b(g5036), .a(n1216) );
  and2_831 AND2_723 ( .c(g10503), .b(g9995), .a(n1337) );
  and2_830 AND2_724 ( .c(g8010), .b(g7738), .a(n1245) );
  and2_829 AND2_725 ( .c(g8410), .b(g713), .a(n1211) );
  and2_828 AND2_726 ( .c(g6231), .b(g818), .a(g5608) );
  and2_827 AND2_727 ( .c(g10581), .b(g10336), .a(n1224) );
  and2_826 AND2_728 ( .c(g10450), .b(g10364), .a(n1071) );
  and2_825 AND2_729 ( .c(g2804), .b(g2132), .a(g1891) );
  and2_824 AND2_730 ( .c(g3418), .b(g2379), .a(g109) );
  and2_823 AND2_731 ( .c(g4820), .b(g186), .a(n1386) );
  and2_822 AND2_732 ( .c(g9653), .b(g1185), .a(g9125) );
  and2_821 AND2_733 ( .c(g6205), .b(g1515), .a(g5151) );
  and2_820 AND2_734 ( .c(g10818), .b(n1225), .a(n1254) );
  and2_819 AND2_735 ( .c(g8172), .b(g37), .a(n1173) );
  and2_818 AND2_736 ( .c(g10496), .b(g10429), .a(n1071) );
  and2_817 AND2_737 ( .c(g5074), .b(g1771), .a(n1202) );
  and2_816 AND2_738 ( .c(g9869), .b(g1558), .a(g9324) );
  and2_815 AND2_739 ( .c(g9719), .b(g1543), .a(n1207) );
  and2_814 AND2_740 ( .c(g10741), .b(g10635), .a(n1365) );
  and2_813 AND2_741 ( .c(g3381), .b(g940), .a(g2756) );
  and2_812 AND2_742 ( .c(g5863), .b(g255), .a(g622) );
  and2_811 AND2_743 ( .c(g8693), .b(n1280), .a(n1174) );
  and2_810 AND2_744 ( .c(g5480), .b(g554), .a(n1389) );
  and2_809 AND2_745 ( .c(g4581), .b(g3766), .a(n1084) );
  and2_808 AND2_746 ( .c(g3685), .b(n1339), .a(g2981) );
  and2_807 AND2_747 ( .c(g5569), .b(g4816), .a(n1150) );
  and2_806 AND2_748 ( .c(g8555), .b(g8409), .a(g7638) );
  and2_805 AND2_749 ( .c(g3263), .b(n1147), .a(n1045) );
  and2_804 AND2_750 ( .c(g9364), .b(g965), .a(n1324) );
  and2_803 AND2_751 ( .c(g4784), .b(g506), .a(g109) );
  and2_802 AND2_752 ( .c(g9454), .b(g8994), .a(g48) );
  and4_11 AND4_5 ( .e(I6331), .d(n1154), .c(n1119), .b(n1118), .a(n1073) );
  and2_801 AND2_753 ( .c(g11299), .b(g4576), .a(n1353) );
  and2_800 AND2_754 ( .c(g6983), .b(g6592), .a(n1083) );
  and2_799 AND2_755 ( .c(g7958), .b(g736), .a(n1251) );
  and2_798 AND2_756 ( .c(g4995), .b(g1474), .a(g4640) );
  and2_797 AND2_757 ( .c(g4079), .b(g1806), .a(g2276) );
  and2_796 AND2_758 ( .c(g2264), .b(g1771), .a(n1333) );
  and2_795 AND2_759 ( .c(g2160), .b(g745), .a(g746) );
  and2_794 AND2_760 ( .c(g3257), .b(g378), .a(g2496) );
  and2_793 AND2_761 ( .c(g3101), .b(I6309), .a(I6310) );
  and2_792 AND2_762 ( .c(g5000), .b(g1470), .a(g4640) );
  and2_791 AND2_763 ( .c(g3301), .b(g1346), .a(g2544) );
  and2_790 AND2_764 ( .c(g5126), .b(g1104), .a(n1235) );
  and4_10 AND4_6 ( .e(I5084), .d(g1462), .c(g1470), .b(g1474), .a(g1478) );
  and2_789 AND2_765 ( .c(g9412), .b(g1727), .a(g9052) );
  and2_788 AND2_766 ( .c(g9389), .b(g1330), .a(n1325) );
  and2_787 AND2_767 ( .c(g2379), .b(g744), .a(g743) );
  and2_786 AND2_768 ( .c(g10706), .b(g10567), .a(n1365) );
  and3_22 AND3_27 ( .d(I16145), .c(g10366), .b(g10447), .a(g10446) );
  and2_785 AND2_769 ( .c(g10597), .b(g10533), .a(n1159) );
  and3_21 AND3_28 ( .d(g8965), .c(n1283), .b(n1307), .a(n1274) );
  and2_784 AND2_770 ( .c(g5608), .b(g814), .a(g4831) );
  and2_783 AND2_771 ( .c(g5220), .b(g1083), .a(n1161) );
  and2_782 AND2_772 ( .c(g10624), .b(g10494), .a(n1159) );
  and2_781 AND2_773 ( .c(g10300), .b(n1224), .a(g10019) );
  and2_780 AND2_774 ( .c(g5023), .b(g1071), .a(n1161) );
  and2_779 AND2_775 ( .c(g4432), .b(n1279), .a(n1055) );
  and2_778 AND2_776 ( .c(g4053), .b(g1786), .a(g2276) );
  and2_777 AND2_777 ( .c(g8050), .b(g7596), .a(g5919) );
  and2_776 AND2_778 ( .c(g5588), .b(g1639), .a(n1389) );
  and3_20 AND3_29 ( .d(g6679), .c(n1295), .b(g6074), .a(g109) );
  and2_775 AND2_779 ( .c(g9963), .b(g9953), .a(n1319) );
  and2_774 AND2_780 ( .c(g3772), .b(n1069), .a(g3089) );
  and2_773 AND2_781 ( .c(g5051), .b(g4432), .a(n1128) );
  and2_772 AND2_782 ( .c(g6831), .b(g207), .a(g5354) );
  and2_771 AND2_783 ( .c(g2981), .b(g1776), .a(g2264) );
  and2_770 AND2_784 ( .c(g8724), .b(g8214), .a(n1384) );
  and2_769 AND2_785 ( .c(g4157), .b(g1796), .a(n1103) );
  and2_768 AND2_786 ( .c(g9707), .b(g1583), .a(n1190) );
  and3_19 AND3_30 ( .d(g8878), .c(n1242), .b(n1307), .a(n1281) );
  and2_767 AND2_787 ( .c(g2132), .b(g1872), .a(g1882) );
  and2_766 AND2_788 ( .c(g10763), .b(g10639), .a(n1365) );
  and3_18 AND3_31 ( .d(g8289), .c(g6777), .b(g8109), .a(n1307) );
  and2_765 AND2_789 ( .c(g7898), .b(g7511), .a(n1253) );
  and2_764 AND2_790 ( .c(g11271), .b(g4753), .a(n1353) );
  and2_763 AND2_791 ( .c(g11461), .b(g11225), .a(g4421) );
  and2_762 AND2_792 ( .c(g5732), .b(g1604), .a(n1215) );
  and2_761 AND2_793 ( .c(g11145), .b(g315), .a(n1354) );
  and2_760 AND2_794 ( .c(g11031), .b(g411), .a(n1347) );
  and2_759 AND2_795 ( .c(g9865), .b(g1607), .a(g9331) );
  and2_758 AND2_796 ( .c(g5944), .b(g1796), .a(g5233) );
  and2_757 AND2_797 ( .c(g9715), .b(g1531), .a(n1207) );
  and2_756 AND2_798 ( .c(g9604), .b(g1194), .a(g9111) );
  and2_755 AND2_799 ( .c(g8799), .b(g8647), .a(n1213) );
  and2_754 AND2_800 ( .c(g11198), .b(g4778), .a(n1354) );
  and2_753 AND2_801 ( .c(g6873), .b(g3263), .a(n1267) );
  and2_752 AND2_802 ( .c(g6632), .b(g61), .a(n1176) );
  and2_751 AND2_803 ( .c(g6095), .b(g1062), .a(g85) );
  and2_750 AND2_804 ( .c(g3863), .b(g1703), .a(g1696) );
  and2_749 AND2_805 ( .c(g9833), .b(g9729), .a(g9785) );
  and2_748 AND2_806 ( .c(g6653), .b(g70), .a(n1176) );
  and2_747 AND2_807 ( .c(g6102), .b(g1038), .a(g85) );
  and2_746 AND2_808 ( .c(g7819), .b(g1887), .a(n1257) );
  and2_745 AND2_809 ( .c(g11393), .b(g11280), .a(n1237) );
  and2_744 AND2_810 ( .c(g2511), .b(n1332), .a(n1336) );
  and2_743 AND2_811 ( .c(g7088), .b(n1137), .a(n1276) );
  and2_742 AND2_812 ( .c(g9584), .b(g1341), .a(n1328) );
  and2_741 AND2_813 ( .c(g9896), .b(g9696), .a(g9624) );
  and3_17 AND3_32 ( .d(g8209), .c(n1222), .b(n1285), .a(n1248) );
  and2_740 AND2_814 ( .c(g6752), .b(g6187), .a(n1056) );
  and2_739 AND2_815 ( .c(g4778), .b(g421), .a(g109) );
  and2_738 AND2_816 ( .c(g11161), .b(n1100), .a(g10937) );
  and2_737 AND2_817 ( .c(g9268), .b(n1385), .a(g8947) );
  and2_736 AND2_818 ( .c(g5681), .b(g135), .a(g5361) );
  and2_735 AND2_819 ( .c(g7951), .b(g73), .a(n1383) );
  and2_734 AND2_820 ( .c(g9419), .b(g1744), .a(n1329) );
  and2_733 AND2_821 ( .c(g10268), .b(n1218), .a(g109) );
  and2_732 AND2_822 ( .c(g5533), .b(g1724), .a(n1185) );
  and2_731 AND2_823 ( .c(g9052), .b(g8936), .a(g48) );
  and2_730 AND2_824 ( .c(g6786), .b(g178), .a(g5919) );
  and2_729 AND2_825 ( .c(g10670), .b(g10396), .a(g8574) );
  and2_728 AND2_826 ( .c(g11087), .b(g829), .a(g10950) );
  and2_727 AND2_827 ( .c(g4949), .b(n1094), .a(n1277) );
  and2_726 AND2_828 ( .c(g6364), .b(g5851), .a(n1365) );
  and2_725 AND2_829 ( .c(g7825), .b(g1941), .a(n1257) );
  and2_724 AND2_830 ( .c(g3400), .b(g115), .a(n1386) );
  and2_723 AND2_831 ( .c(g4998), .b(g1304), .a(g109) );
  and2_722 AND2_832 ( .c(g10667), .b(g10405), .a(n1224) );
  and2_721 AND2_833 ( .c(g7136), .b(g5190), .a(n1199) );
  and2_720 AND2_834 ( .c(g6532), .b(g339), .a(n1176) );
  and2_719 AND2_835 ( .c(g9385), .b(g1324), .a(n1325) );
  and4_9 AND4_7 ( .e(I5690), .d(g1436), .c(g1440), .b(g1444), .a(g1448) );
  and2_718 AND2_836 ( .c(g4484), .b(g1137), .a(g109) );
  and2_717 AND2_837 ( .c(g9897), .b(g9699), .a(g9624) );
  and2_716 AND2_838 ( .c(g9425), .b(g1753), .a(n1329) );
  and2_715 AND2_839 ( .c(g3383), .b(g186), .a(n1386) );
  and2_714 AND2_840 ( .c(g5601), .b(g1035), .a(n1378) );
  and2_713 AND2_841 ( .c(g7943), .b(g64), .a(n1383) );
  and2_712 AND2_842 ( .c(g11171), .b(g481), .a(n1347) );
  and2_711 AND2_843 ( .c(g3423), .b(I6630), .a(I6631) );
  and2_710 AND2_844 ( .c(g7230), .b(g6064), .a(n1276) );
  and2_709 AND2_845 ( .c(g4952), .b(g1648), .a(n1202) );
  and2_708 AND2_846 ( .c(g8736), .b(n1231), .a(g8451) );
  and2_707 AND2_847 ( .c(g6787), .b(g266), .a(n1221) );
  and3_16 AND3_33 ( .d(g8968), .c(n1268), .b(n1307), .a(n1274) );
  and2_706 AND2_848 ( .c(g10306), .b(g10007), .a(g8574) );
  and2_705 AND2_849 ( .c(g9331), .b(g8972), .a(g48) );
  and2_704 AND2_850 ( .c(g11459), .b(g11221), .a(g4421) );
  and2_703 AND2_851 ( .c(g4561), .b(g538), .a(g109) );
  and2_702 AND2_852 ( .c(g11425), .b(g10583), .a(n1200) );
  and2_701 AND2_853 ( .c(g11458), .b(g11219), .a(g4421) );
  and2_700 AND2_854 ( .c(g5739), .b(g1607), .a(n1215) );
  and2_699 AND2_855 ( .c(g7496), .b(n1384), .a(g64) );
  and2_698 AND2_856 ( .c(g4986), .b(g1411), .a(g4682) );
  and2_697 AND2_857 ( .c(g11010), .b(g5187), .a(n1347) );
  and2_696 AND2_858 ( .c(g3999), .b(g1741), .a(n1206) );
  and2_695 AND2_859 ( .c(g8175), .b(g39), .a(n1173) );
  and2_694 AND2_860 ( .c(g8722), .b(g8210), .a(n1384) );
  and2_693 AND2_861 ( .c(g4764), .b(g411), .a(g109) );
  and2_692 AND2_862 ( .c(g7137), .b(g5590), .a(n1236) );
  and2_691 AND2_863 ( .c(g7891), .b(g7471), .a(n1253) );
  and2_690 AND2_864 ( .c(g8651), .b(g8261), .a(n1365) );
  and2_689 AND2_865 ( .c(g5479), .b(g1845), .a(n1288) );
  and2_688 AND2_866 ( .c(g11599), .b(g1341), .a(n1192) );
  and2_687 AND2_867 ( .c(g6684), .b(g91), .a(n1316) );
  and2_686 AND2_868 ( .c(g6745), .b(g5605), .a(g5557) );
  and2_685 AND2_869 ( .c(g6639), .b(g357), .a(n1176) );
  and2_684 AND2_870 ( .c(g10937), .b(n1172), .a(n1347) );
  and2_683 AND2_871 ( .c(g3696), .b(g1713), .a(n1364) );
  and2_682 AND2_872 ( .c(g4503), .b(g654), .a(n1089) );
  and2_681 AND2_873 ( .c(g6791), .b(g269), .a(n1221) );
  and2_680 AND2_874 ( .c(g5190), .b(g1245), .a(g109) );
  and2_679 AND2_875 ( .c(g5390), .b(g1101), .a(n1235) );
  and2_678 AND2_876 ( .c(g8384), .b(g8180), .a(n1386) );
  and2_677 AND2_877 ( .c(g4224), .b(g1092), .a(n1364) );
  and2_676 AND2_878 ( .c(g5501), .b(g1672), .a(n1378) );
  and2_675 AND2_879 ( .c(g9173), .b(g8968), .a(g48) );
  and2_674 AND2_880 ( .c(g6759), .b(g148), .a(g5919) );
  and2_673 AND2_881 ( .c(g8838), .b(g8602), .a(n1233) );
  and2_672 AND2_882 ( .c(g8024), .b(g6577), .a(n1277) );
  and2_671 AND2_883 ( .c(g10666), .b(g10402), .a(n1224) );
  and2_670 AND2_884 ( .c(g11158), .b(g309), .a(n1354) );
  and2_669 AND2_885 ( .c(g9602), .b(g932), .a(n1326) );
  and2_668 AND2_886 ( .c(g5704), .b(g143), .a(g5361) );
  and2_667 AND2_887 ( .c(g4617), .b(g3275), .a(g3879) );
  and2_666 AND2_888 ( .c(g11561), .b(g11492), .a(n1364) );
  and2_665 AND2_889 ( .c(g9868), .b(g1555), .a(g9324) );
  and2_664 AND2_890 ( .c(g11295), .b(g4554), .a(n1354) );
  and2_663 AND2_891 ( .c(g11144), .b(g305), .a(n1357) );
  and2_662 AND2_892 ( .c(g9718), .b(g1540), .a(n1207) );
  and2_661 AND2_893 ( .c(g3434), .b(g237), .a(n1386) );
  and2_660 AND2_894 ( .c(g4987), .b(g1440), .a(g4682) );
  and2_659 AND2_895 ( .c(g4771), .b(g496), .a(g109) );
  and2_658 AND2_896 ( .c(g5250), .b(g1270), .a(g109) );
  and2_657 AND2_897 ( .c(g6098), .b(g1065), .a(g85) );
  and2_656 AND2_898 ( .c(g9582), .b(g1336), .a(n1328) );
  and2_655 AND2_899 ( .c(g6833), .b(g186), .a(g5354) );
  and2_654 AND2_900 ( .c(g3533), .b(n1140), .a(g2892) );
  and2_653 AND2_901 ( .c(g4892), .b(g632), .a(n1263) );
  and2_652 AND2_902 ( .c(g8104), .b(g5493), .a(g6740) );
  and2_651 AND2_903 ( .c(g9415), .b(g1733), .a(g9052) );
  and2_650 AND2_904 ( .c(g8499), .b(g8377), .a(g3041) );
  and2_649 AND2_905 ( .c(g9664), .b(g1191), .a(g9125) );
  and2_648 AND2_906 ( .c(g10740), .b(n1294), .a(n1298) );
  and2_647 AND2_907 ( .c(g2534), .b(g798), .a(g794) );
  and2_646 AND2_908 ( .c(g8754), .b(n1231), .a(g8451) );
  and2_645 AND2_909 ( .c(g9721), .b(g9413), .a(n1386) );
  and2_644 AND2_910 ( .c(g6162), .b(g3584), .a(g3374) );
  and2_643 AND2_911 ( .c(g4991), .b(g1508), .a(g4640) );
  and2_642 AND2_912 ( .c(g6362), .b(g5846), .a(n1364) );
  and4_8 AND4_8 ( .e(I6631), .d(g1791), .c(g1796), .b(g1801), .a(g1806) );
  and2_641 AND2_913 ( .c(g10685), .b(g10383), .a(g3863) );
  and2_640 AND2_914 ( .c(g4340), .b(g1153), .a(g109) );
  and2_639 AND2_915 ( .c(g11023), .b(g440), .a(n1348) );
  and2_638 AND2_916 ( .c(g8044), .b(g7598), .a(g5919) );
  and2_637 AND2_917 ( .c(g11224), .b(g968), .a(n1177) );
  and2_636 AND2_918 ( .c(g11571), .b(n1123), .a(g11561) );
  and2_635 AND2_919 ( .c(g4959), .b(g1520), .a(g4682) );
  and2_634 AND2_920 ( .c(g10334), .b(n1217), .a(g109) );
  and2_633 AND2_921 ( .c(g5626), .b(g1633), .a(n1391) );
  and2_632 AND2_922 ( .c(g9940), .b(g9920), .a(n1320) );
  and2_631 AND2_923 ( .c(g4876), .b(g1086), .a(n1364) );
  and2_630 AND2_924 ( .c(g6728), .b(g4482), .a(n1286) );
  and2_629 AND2_925 ( .c(g6730), .b(g1872), .a(g5013) );
  and2_628 AND2_926 ( .c(g9689), .b(g263), .a(n1171) );
  and2_627 AND2_927 ( .c(g10762), .b(g10635), .a(n1364) );
  and2_626 AND2_928 ( .c(g6070), .b(g1050), .a(g85) );
  and2_625 AND2_929 ( .c(g9428), .b(g1756), .a(n1329) );
  and2_624 AND2_930 ( .c(g9030), .b(g8935), .a(g48) );
  and2_623 AND2_931 ( .c(g9430), .b(g1759), .a(n1329) );
  and2_622 AND2_932 ( .c(g8927), .b(n1307), .a(g8642) );
  and2_621 AND2_933 ( .c(g7068), .b(g5024), .a(n1199) );
  and2_620 AND2_934 ( .c(g8014), .b(g7740), .a(n1245) );
  and2_619 AND2_935 ( .c(g11392), .b(g11278), .a(n1237) );
  and2_618 AND2_936 ( .c(g5782), .b(g1558), .a(n1229) );
  and2_617 AND2_937 ( .c(g9910), .b(n1182), .a(n1327) );
  and2_616 AND2_938 ( .c(g4824), .b(g774), .a(g4099) );
  and2_615 AND2_939 ( .c(g6331), .b(g201), .a(g5354) );
  and2_614 AND2_940 ( .c(g4236), .b(g1098), .a(n1364) );
  and2_613 AND2_941 ( .c(g11559), .b(g1801), .a(g11519) );
  and2_612 AND2_942 ( .c(g9609), .b(g907), .a(g9205) );
  and2_611 AND2_943 ( .c(g11558), .b(g1796), .a(g11519) );
  and2_610 AND2_944 ( .c(g6087), .b(g1056), .a(g85) );
  and2_609 AND2_945 ( .c(g4877), .b(g243), .a(n1386) );
  and2_608 AND2_946 ( .c(g5526), .b(g1950), .a(g3209) );
  and2_607 AND2_947 ( .c(g10751), .b(g10646), .a(n1364) );
  and2_606 AND2_948 ( .c(g10772), .b(g10655), .a(n1364) );
  and2_605 AND2_949 ( .c(g8135), .b(g1945), .a(n1210) );
  and2_604 AND2_950 ( .c(g11544), .b(n1293), .a(n1299) );
  and2_603 AND2_951 ( .c(g5084), .b(g1776), .a(n1202) );
  and2_602 AND2_952 ( .c(g8382), .b(g5248), .a(g7101) );
  and2_601 AND2_953 ( .c(g10230), .b(n1224), .a(g9968) );
  and2_600 AND2_954 ( .c(g5484), .b(g1896), .a(g3209) );
  and2_599 AND2_955 ( .c(g7241), .b(g6772), .a(g5557) );
  and2_598 AND2_956 ( .c(g3942), .b(g219), .a(g2355) );
  and2_597 AND2_957 ( .c(g10638), .b(g10383), .a(g3829) );
  and2_596 AND2_958 ( .c(g4064), .b(g1759), .a(n1206) );
  and2_595 AND2_959 ( .c(g9365), .b(g1321), .a(n1325) );
  and2_594 AND2_960 ( .c(g9861), .b(g9738), .a(g9579) );
  and2_593 AND2_961 ( .c(g8749), .b(n1234), .a(g8488) );
  and2_592 AND2_962 ( .c(g11255), .b(n1336), .a(n1191) );
  and2_591 AND2_963 ( .c(g11189), .b(g4736), .a(n1357) );
  and2_590 AND2_964 ( .c(g10510), .b(g10019), .a(n1337) );
  and3_15 AND3_34 ( .d(g8947), .c(n1247), .b(n1307), .a(n1266) );
  and2_589 AND2_965 ( .c(g2917), .b(n1103), .a(g1657) );
  and2_588 AND2_966 ( .c(g5919), .b(n1295), .a(g109) );
  and2_587 AND2_967 ( .c(g11188), .b(g4732), .a(n1355) );
  and2_586 AND2_968 ( .c(g9846), .b(g287), .a(g9313) );
  and2_585 AND2_969 ( .c(g7818), .b(g1878), .a(n1257) );
  and2_584 AND2_970 ( .c(g11460), .b(g11223), .a(g4421) );
  and2_583 AND2_971 ( .c(g5276), .b(g736), .a(g3041) );
  and2_582 AND2_972 ( .c(g11030), .b(g406), .a(n1348) );
  and2_581 AND2_973 ( .c(g11093), .b(g841), .a(g10950) );
  and2_580 AND2_974 ( .c(g7893), .b(g7478), .a(n1253) );
  and2_579 AND2_975 ( .c(g8653), .b(g8265), .a(n1364) );
  and2_578 AND2_976 ( .c(g10442), .b(g9968), .a(n1337) );
  and2_577 AND2_977 ( .c(g6535), .b(g345), .a(n1176) );
  and2_576 AND2_978 ( .c(g8102), .b(g5485), .a(g6740) );
  and4_7 AND4_9 ( .e(I5085), .d(g1490), .c(g1494), .b(g1504), .a(g1508) );
  and2_575 AND2_979 ( .c(g5004), .b(g1296), .a(g109) );
  and2_574 AND2_980 ( .c(g3912), .b(g207), .a(g2355) );
  and2_573 AND2_981 ( .c(g7186), .b(n1147), .a(n1267) );
  and2_572 AND2_982 ( .c(g4489), .b(g348), .a(g3586) );
  and2_571 AND2_983 ( .c(g9662), .b(g123), .a(n1331) );
  and2_570 AND2_984 ( .c(g9418), .b(g1741), .a(g9052) );
  and2_569 AND2_985 ( .c(g11218), .b(g959), .a(n1177) );
  and2_568 AND2_986 ( .c(g4471), .b(g1121), .a(g109) );
  and2_567 AND2_987 ( .c(g10746), .b(g10643), .a(n1364) );
  and2_566 AND2_988 ( .c(g7125), .b(g1212), .a(g5763) );
  and2_565 AND2_989 ( .c(g7821), .b(g1905), .a(n1257) );
  and2_564 AND2_990 ( .c(g6246), .b(g178), .a(g5361) );
  and2_563 AND2_991 ( .c(g9256), .b(n1385), .a(g8963) );
  and2_562 AND2_992 ( .c(g8042), .b(g7533), .a(g5128) );
  and2_561 AND2_993 ( .c(g10237), .b(g9968), .a(g8574) );
  and2_560 AND2_994 ( .c(g7939), .b(g61), .a(n1383) );
  and2_559 AND2_995 ( .c(g8786), .b(g8638), .a(n1213) );
  and2_558 AND2_996 ( .c(g10684), .b(g10382), .a(g3863) );
  and2_557 AND2_997 ( .c(g11455), .b(g11233), .a(g4421) );
  and2_556 AND2_998 ( .c(g8364), .b(g658), .a(n1211) );
  and3_14 AND3_35 ( .d(g2990), .c(n1131), .b(n1093), .a(g1814) );
  and2_555 AND2_999 ( .c(g9847), .b(g290), .a(g9313) );
  and2_554 AND2_1000 ( .c(g8054), .b(g7584), .a(g5919) );
  and2_553 AND2_1001 ( .c(g5617), .b(g1050), .a(n1378) );
  and2_552 AND2_1002 ( .c(g6502), .b(g5981), .a(n1083) );
  and2_551 AND2_1003 ( .c(g5789), .b(g1561), .a(n1229) );
  and2_550 AND2_1004 ( .c(g4009), .b(g1747), .a(n1206) );
  and2_549 AND2_1005 ( .c(g11277), .b(g4779), .a(n1352) );
  and2_548 AND2_1006 ( .c(g6940), .b(g6472), .a(g1945) );
  and2_547 AND2_1007 ( .c(g7061), .b(g790), .a(g6760) );
  and2_546 AND2_1008 ( .c(g11595), .b(g1336), .a(n1192) );
  and2_545 AND2_1009 ( .c(g5771), .b(g1534), .a(n1229) );
  and2_544 AND2_1010 ( .c(g8553), .b(g8405), .a(g7638) );
  and2_543 AND2_1011 ( .c(g4836), .b(g643), .a(n1089) );
  and2_542 AND2_1012 ( .c(g5547), .b(g1733), .a(n1185) );
  and2_541 AND2_1013 ( .c(g6216), .b(g1407), .a(g5151) );
  and2_540 AND2_1014 ( .c(g4967), .b(g1515), .a(g4682) );
  and2_539 AND2_1015 ( .c(g6671), .b(g342), .a(n1176) );
  and2_538 AND2_1016 ( .c(g7200), .b(g3098), .a(n1276) );
  and2_537 AND2_1017 ( .c(g3661), .b(g382), .a(g3257) );
  and2_536 AND2_1018 ( .c(g7046), .b(g4998), .a(n1199) );
  and2_535 AND2_1019 ( .c(g4229), .b(g999), .a(n1378) );
  and2_534 AND2_1020 ( .c(g8389), .b(g5263), .a(g7101) );
  and2_533 AND2_1021 ( .c(g6430), .b(g5044), .a(g5013) );
  and2_532 AND2_1022 ( .c(g8706), .b(n1234), .a(g8488) );
  and2_531 AND2_1023 ( .c(g4993), .b(g1448), .a(g4682) );
  and2_530 AND2_1024 ( .c(g6247), .b(g127), .a(g5361) );
  and2_529 AND2_1025 ( .c(g9257), .b(n1385), .a(g8964) );
  and2_528 AND2_1026 ( .c(g11170), .b(g525), .a(n1348) );
  and2_527 AND2_1027 ( .c(g7145), .b(g5250), .a(n1199) );
  and2_526 AND2_1028 ( .c(g5738), .b(g1586), .a(n1215) );
  and2_525 AND2_1029 ( .c(g6826), .b(g225), .a(g5354) );
  and2_524 AND2_1030 ( .c(g7191), .b(g5219), .a(n1286) );
  and2_523 AND2_1031 ( .c(g3998), .b(n1333), .a(g2276) );
  and2_522 AND2_1032 ( .c(g6741), .b(g3284), .a(g5557) );
  and2_521 AND2_1033 ( .c(g5478), .b(g1905), .a(g3209) );
  and2_520 AND2_1034 ( .c(g11167), .b(g538), .a(n1348) );
  and2_519 AND2_1035 ( .c(g11194), .b(g4764), .a(n1355) );
  and2_518 AND2_1036 ( .c(g11589), .b(g1333), .a(n1198) );
  and2_517 AND2_1037 ( .c(g6638), .b(g64), .a(n1176) );
  and2_516 AND2_1038 ( .c(g4921), .b(g627), .a(g4431) );
  and2_515 AND2_1039 ( .c(g7536), .b(n1384), .a(g76) );
  and2_514 AND2_1040 ( .c(g9585), .b(g889), .a(g8995) );
  and2_513 AND2_1041 ( .c(g2957), .b(n1103), .a(g1663) );
  and2_512 AND2_1042 ( .c(g11588), .b(g1330), .a(n1198) );
  and2_511 AND2_1043 ( .c(g5690), .b(g1567), .a(n1215) );
  and2_510 AND2_1044 ( .c(g6883), .b(g1923), .a(g6003) );
  and2_509 AND2_1045 ( .c(g4837), .b(g1068), .a(n1364) );
  and3_13 AND3_36 ( .d(g8963), .c(n1247), .b(n1307), .a(n1274) );
  and2_508 AND2_1046 ( .c(g8791), .b(g8641), .a(n1213) );
  and2_507 AND2_1047 ( .c(g6217), .b(g563), .a(n1379) );
  and4_6 AND4_10 ( .e(I6316), .d(n1061), .c(n1074), .b(n1082), .a(n1086) );
  and2_506 AND2_1048 ( .c(g11022), .b(g444), .a(n1348) );
  and2_505 AND2_1049 ( .c(g5915), .b(g4168), .a(g4977) );
  and2_504 AND2_1050 ( .c(g4788), .b(g511), .a(g109) );
  and2_503 AND2_1051 ( .c(g8759), .b(n1231), .a(g8451) );
  and2_502 AND2_1052 ( .c(g5110), .b(g1806), .a(n1202) );
  and2_501 AND2_1053 ( .c(g11254), .b(g986), .a(n1169) );
  and2_500 AND2_1054 ( .c(g6827), .b(g219), .a(g5354) );
  and3_12 AND3_37 ( .d(g8957), .c(n1284), .b(n1307), .a(n1266) );
  and2_499 AND2_1055 ( .c(g6333), .b(g197), .a(g5354) );
  and2_498 AND2_1056 ( .c(g8049), .b(g7567), .a(g5919) );
  and2_497 AND2_1057 ( .c(g4392), .b(g3273), .a(g3829) );
  and2_496 AND2_1058 ( .c(g9856), .b(g1592), .a(g9331) );
  and2_495 AND2_1059 ( .c(g9411), .b(g1724), .a(g9052) );
  and2_494 AND2_1060 ( .c(g5002), .b(g1494), .a(g4640) );
  and2_493 AND2_1061 ( .c(g11101), .b(g857), .a(g10950) );
  and2_492 AND2_1062 ( .c(g11177), .b(g511), .a(n1348) );
  and2_491 AND2_1063 ( .c(g11560), .b(g1806), .a(g11519) );
  and2_490 AND2_1064 ( .c(g8098), .b(g5478), .a(g6740) );
  and2_489 AND2_1065 ( .c(g3970), .b(g225), .a(g2355) );
  and2_488 AND2_1066 ( .c(g4941), .b(g1038), .a(n1379) );
  and2_487 AND2_1067 ( .c(g10453), .b(n1166), .a(n1071) );
  and2_486 AND2_1068 ( .c(g5877), .b(g4921), .a(g639) );
  and2_485 AND2_1069 ( .c(g6662), .b(g366), .a(n1176) );
  and2_484 AND2_1070 ( .c(g7935), .b(g58), .a(n1383) );
  and2_483 AND2_1071 ( .c(g6067), .b(g1047), .a(g85) );
  and4_5 AND4_11 ( .e(I6317), .d(n1077), .c(n1113), .b(n1065), .a(n1053) );
  and2_482 AND2_1072 ( .c(g9863), .b(g9740), .a(g9052) );
  and4_4 AND4_12 ( .e(I5886), .d(g174), .c(g170), .b(n1156), .a(n1146) );
  and2_481 AND2_1073 ( .c(g6994), .b(g6758), .a(g3829) );
  and2_480 AND2_1074 ( .c(g9713), .b(g1589), .a(n1190) );
  and2_479 AND2_1075 ( .c(g4431), .b(n1091), .a(g3533) );
  and2_478 AND2_1076 ( .c(g4252), .b(g1007), .a(n1379) );
  and2_477 AND2_1077 ( .c(g11166), .b(g542), .a(n1348) );
  and2_476 AND2_1078 ( .c(g7130), .b(g5150), .a(n1199) );
  and2_475 AND2_1079 ( .c(g11009), .b(g5179), .a(n1348) );
  and2_474 AND2_1080 ( .c(g7542), .b(n1384), .a(g79) );
  and2_473 AND2_1081 ( .c(g8019), .b(g6573), .a(n1286) );
  and2_472 AND2_1082 ( .c(g11008), .b(g5171), .a(n1348) );
  and2_471 AND2_1083 ( .c(g3516), .b(g1209), .a(n1363) );
  and2_470 AND2_1084 ( .c(g8052), .b(g7573), .a(g5128) );
  and2_469 AND2_1085 ( .c(g3987), .b(g243), .a(g2355) );
  and2_468 AND2_1086 ( .c(g4765), .b(g491), .a(g109) );
  and2_467 AND2_1087 ( .c(g11555), .b(n1339), .a(g11519) );
  and2_466 AND2_1088 ( .c(g9857), .b(g9734), .a(g9569) );
  and2_465 AND2_1089 ( .c(g8728), .b(g8226), .a(n1384) );
  and2_464 AND2_1090 ( .c(g8730), .b(g8230), .a(n1384) );
  and2_463 AND2_1091 ( .c(g8185), .b(g664), .a(g7101) );
  and2_462 AND2_1092 ( .c(g5194), .b(g1610), .a(n1202) );
  and2_461 AND2_1093 ( .c(g8385), .b(g5255), .a(g7101) );
  and2_460 AND2_1094 ( .c(g4610), .b(g3804), .a(n1117) );
  and2_459 AND2_1095 ( .c(g7902), .b(g7661), .a(n1276) );
  and2_458 AND2_1096 ( .c(g4073), .b(g3200), .a(g3222) );
  and2_457 AND2_1097 ( .c(g8070), .b(g682), .a(n1251) );
  and2_456 AND2_1098 ( .c(g5731), .b(g1583), .a(n1215) );
  and2_455 AND2_1099 ( .c(g11238), .b(g4553), .a(n1355) );
  and2_454 AND2_1100 ( .c(g4473), .b(g1125), .a(g109) );
  and2_453 AND2_1101 ( .c(g8470), .b(g8308), .a(g7246) );
  and2_452 AND2_1102 ( .c(g5489), .b(g557), .a(n1391) );
  and2_451 AND2_1103 ( .c(g3991), .b(g1738), .a(n1206) );
  and4_3 AND4_13 ( .e(I5887), .d(n1152), .c(n1136), .b(g166), .a(n1108) );
  and2_450 AND2_1104 ( .c(g7823), .b(g1923), .a(n1257) );
  and2_449 AND2_1105 ( .c(g4069), .b(g1762), .a(n1206) );
  and3_11 AND3_38 ( .d(g11519), .c(g1317), .b(n1367), .a(g11492) );
  and2_448 AND2_1106 ( .c(g11176), .b(g506), .a(n1348) );
  and2_447 AND2_1107 ( .c(g11092), .b(g837), .a(g10950) );
  and2_446 AND2_1108 ( .c(g11154), .b(g330), .a(n1355) );
  and2_445 AND2_1109 ( .c(g9608), .b(g7), .a(n1331) );
  and2_444 AND2_1110 ( .c(g11637), .b(n1212), .a(g4421) );
  and2_443 AND2_1111 ( .c(g2091), .b(g976), .a(g971) );
  and2_442 AND2_1112 ( .c(g8406), .b(g695), .a(n1211) );
  and2_441 AND2_1113 ( .c(g5254), .b(g549), .a(n1391) );
  and2_440 AND2_1114 ( .c(g7260), .b(g6752), .a(n1092) );
  and2_439 AND2_1115 ( .c(g5150), .b(g1275), .a(g109) );
  and2_438 AND2_1116 ( .c(g8766), .b(g8612), .a(g5151) );
  and2_437 AND2_1117 ( .c(g9588), .b(g1351), .a(n1328) );
  and2_436 AND2_1118 ( .c(g8801), .b(g8742), .a(n1213) );
  and2_435 AND2_1119 ( .c(g7063), .b(g5008), .a(n1199) );
  and2_434 AND2_1120 ( .c(g10303), .b(g9995), .a(g8574) );
  and2_433 AND2_1121 ( .c(g5009), .b(g1486), .a(g4640) );
  and2_432 AND2_1122 ( .c(g9665), .b(g1314), .a(n1325) );
  and2_431 AND2_1123 ( .c(g8748), .b(n1234), .a(g8488) );
  and2_430 AND2_1124 ( .c(g11215), .b(g953), .a(n1177) );
  and2_429 AND2_1125 ( .c(g10750), .b(g10597), .a(g3586) );
  and3_10 AND3_39 ( .d(g5769), .c(n1062), .b(g4921), .a(g3818) );
  and2_428 AND2_1126 ( .c(g8755), .b(n1231), .a(g8451) );
  and2_427 AND2_1127 ( .c(g6673), .b(g90), .a(n1316) );
  and2_426 AND2_1128 ( .c(g5212), .b(g1255), .a(g109) );
  and2_425 AND2_1129 ( .c(g7720), .b(g727), .a(g6488) );
  and3_9 AND3_40 ( .d(g5918), .c(g109), .b(n1295), .a(g4609) );
  and2_424 AND2_1130 ( .c(g8045), .b(g7547), .a(g5128) );
  and2_423 AND2_1131 ( .c(g8173), .b(g7971), .a(n1083) );
  and2_422 AND2_1132 ( .c(g11349), .b(g11288), .a(n1237) );
  and2_421 AND2_1133 ( .c(g7843), .b(g7599), .a(g5919) );
  and2_420 AND2_1134 ( .c(g9696), .b(g281), .a(n1171) );
  and2_419 AND2_1135 ( .c(g6772), .b(g6228), .a(g722) );
  and2_418 AND2_1136 ( .c(g6058), .b(g1035), .a(g85) );
  and2_417 AND2_1137 ( .c(g6531), .b(g79), .a(n1176) );
  and2_416 AND2_1138 ( .c(g6743), .b(g4106), .a(g5557) );
  and2_415 AND2_1139 ( .c(g6890), .b(g6752), .a(n1267) );
  and2_414 AND2_1140 ( .c(g7549), .b(g7269), .a(g3829) );
  and2_413 AND2_1141 ( .c(g8169), .b(g35), .a(n1173) );
  and2_412 AND2_1142 ( .c(g11304), .b(g4585), .a(n1355) );
  and2_411 AND2_1143 ( .c(g9944), .b(g9924), .a(n1321) );
  and2_410 AND2_1144 ( .c(g9240), .b(g48), .a(g8962) );
  and2_409 AND2_1145 ( .c(g8059), .b(g7592), .a(g5919) );
  and2_408 AND2_1146 ( .c(g8718), .b(g8203), .a(n1384) );
  and2_407 AND2_1147 ( .c(g8767), .b(g8616), .a(g5151) );
  and2_406 AND2_1148 ( .c(g9316), .b(g8877), .a(g48) );
  and2_405 AND2_1149 ( .c(g7625), .b(g673), .a(g6488) );
  and2_404 AND2_1150 ( .c(g8793), .b(g8644), .a(n1213) );
  and2_403 AND2_1151 ( .c(g2940), .b(n1103), .a(g1654) );
  and2_402 AND2_1152 ( .c(g4114), .b(g1351), .a(g3301) );
  and2_401 AND2_1153 ( .c(g11636), .b(g11624), .a(n1238) );
  and2_400 AND2_1154 ( .c(g10949), .b(g2947), .a(g10809) );
  and2_399 AND2_1155 ( .c(g4870), .b(g237), .a(g2355) );
  and2_398 AND2_1156 ( .c(g3563), .b(g3275), .a(n1158) );
  and2_397 AND2_1157 ( .c(g10948), .b(g2223), .a(g10809) );
  and2_396 AND2_1158 ( .c(g8246), .b(g7846), .a(n1245) );
  and2_395 AND2_1159 ( .c(g5788), .b(g1540), .a(n1229) );
  and2_394 AND2_1160 ( .c(g4008), .b(g1776), .a(g2276) );
  and2_393 AND2_1161 ( .c(g9596), .b(g928), .a(n1326) );
  and2_392 AND2_1162 ( .c(g5249), .b(g1089), .a(n1161) );
  and2_391 AND2_1163 ( .c(g11585), .b(g1321), .a(n1198) );
  and2_390 AND2_1164 ( .c(g3089), .b(n1050), .a(n1076) );
  and2_389 AND2_1165 ( .c(g4972), .b(g1436), .a(g4682) );
  and2_388 AND2_1166 ( .c(g11554), .b(g1776), .a(g11519) );
  and2_387 AND2_1167 ( .c(g7586), .b(g7096), .a(n1240) );
  and2_386 AND2_1168 ( .c(g10673), .b(g10417), .a(n1224) );
  and3_8 AND3_41 ( .d(g4806), .c(g3215), .b(g3992), .a(g2493) );
  and2_385 AND2_1169 ( .c(g5485), .b(g1914), .a(g3209) );
  and2_384 AND2_1170 ( .c(g9936), .b(g9915), .a(g9624) );
  and2_383 AND2_1171 ( .c(g2910), .b(n1103), .a(g1660) );
  and2_382 AND2_1172 ( .c(g9317), .b(n1385), .a(g8875) );
  and2_381 AND2_1173 ( .c(g10933), .b(g10853), .a(g1854) );
  and2_380 AND2_1174 ( .c(g8388), .b(g8177), .a(g7246) );
  and2_379 AND2_1175 ( .c(g4465), .b(g1117), .a(g109) );
  and2_378 AND2_1176 ( .c(g7141), .b(g5230), .a(n1199) );
  and2_377 AND2_1177 ( .c(g10508), .b(g10013), .a(n1337) );
  and2_376 AND2_1178 ( .c(g4230), .b(g1095), .a(n1363) );
  and2_375 AND2_1179 ( .c(g10634), .b(g10382), .a(g3829) );
  and2_374 AND2_1180 ( .c(g9601), .b(g922), .a(g9192) );
  and2_373 AND2_1181 ( .c(g6126), .b(g3681), .a(n1277) );
  and2_372 AND2_1182 ( .c(g6326), .b(g1250), .a(n1322) );
  and2_371 AND2_1183 ( .c(g7710), .b(g700), .a(g6488) );
  and2_370 AND2_1184 ( .c(g8028), .b(g7375), .a(n1245) );
  and2_369 AND2_1185 ( .c(g6760), .b(g786), .a(g6221) );
  and2_368 AND2_1186 ( .c(g5640), .b(g1059), .a(n1379) );
  and2_367 AND2_1187 ( .c(g5031), .b(g1478), .a(g4640) );
  and2_366 AND2_1188 ( .c(g4550), .b(g342), .a(g3586) );
  and2_365 AND2_1189 ( .c(g7879), .b(g5286), .a(n1390) );
  and2_364 AND2_1190 ( .c(g7962), .b(g7730), .a(n1267) );
  and2_363 AND2_1191 ( .c(g9597), .b(g1170), .a(g9125) );
  and2_362 AND2_1192 ( .c(g10452), .b(n1194), .a(n1071) );
  and2_361 AND2_1193 ( .c(g4891), .b(g631), .a(n1263) );
  and2_360 AND2_1194 ( .c(g5005), .b(g1490), .a(g4640) );
  and2_359 AND2_1195 ( .c(g6423), .b(g4348), .a(g5013) );
  and2_358 AND2_1196 ( .c(g8108), .b(g1891), .a(n1210) );
  and3_7 AND3_42 ( .d(g4807), .c(n1367), .b(g1289), .a(n1083) );
  and2_357 AND2_1197 ( .c(g5911), .b(g3322), .a(g4977) );
  and2_356 AND2_1198 ( .c(g9937), .b(g9916), .a(g9624) );
  and2_355 AND2_1199 ( .c(g9840), .b(g9704), .a(g9747) );
  and2_354 AND2_1200 ( .c(g10780), .b(g10723), .a(n1202) );
  and2_353 AND2_1201 ( .c(g8217), .b(g1872), .a(n1210) );
  and2_352 AND2_1202 ( .c(g11013), .b(g5209), .a(n1348) );
  and2_351 AND2_1203 ( .c(g9390), .b(g1333), .a(n1325) );
  and2_350 AND2_1204 ( .c(g11214), .b(g950), .a(n1177) );
  and2_349 AND2_1205 ( .c(g6327), .b(g1255), .a(n1322) );
  and2_348 AND2_1206 ( .c(g4342), .b(g1149), .a(g109) );
  and2_347 AND2_1207 ( .c(g5796), .b(g1564), .a(n1229) );
  and2_346 AND2_1208 ( .c(g5473), .b(g546), .a(n1390) );
  and2_345 AND2_1209 ( .c(g6346), .b(g5038), .a(n1216) );
  and2_344 AND2_1210 ( .c(g6633), .b(g354), .a(n1176) );
  and2_343 AND2_1211 ( .c(g11005), .b(g5119), .a(n1348) );
  and2_342 AND2_1212 ( .c(g8365), .b(g668), .a(n1211) );
  and2_341 AND2_1213 ( .c(g8048), .b(g7558), .a(g5919) );
  and2_340 AND2_1214 ( .c(g4481), .b(g1713), .a(n1380) );
  and2_339 AND2_1215 ( .c(g4097), .b(n1333), .a(n1103) );
  and2_338 AND2_1216 ( .c(g8055), .b(g7588), .a(g5128) );
  and2_337 AND2_1217 ( .c(g4497), .b(g351), .a(g3586) );
  and2_336 AND2_1218 ( .c(g9942), .b(g9922), .a(n1320) );
  and2_335 AND2_1219 ( .c(g6696), .b(g94), .a(n1316) );
  and3_6 AND3_43 ( .d(g10731), .c(g5118), .b(g1850), .a(g10665) );
  and2_334 AND2_1220 ( .c(g8827), .b(g8552), .a(n1213) );
  and2_333 AND2_1221 ( .c(g5540), .b(g1727), .a(n1185) );
  and2_332 AND2_1222 ( .c(g4960), .b(g1403), .a(g4682) );
  and2_331 AND2_1223 ( .c(g8846), .b(g8615), .a(n1233) );
  and2_330 AND2_1224 ( .c(g6508), .b(g5983), .a(n1083) );
  and2_329 AND2_1225 ( .c(g6240), .b(g182), .a(g5361) );
  and2_328 AND2_1226 ( .c(g7931), .b(g52), .a(n1383) );
  and2_327 AND2_1227 ( .c(g5287), .b(n1301), .a(n1227) );
  and2_326 AND2_1228 ( .c(g6472), .b(g5853), .a(g1936) );
  and2_325 AND2_1229 ( .c(g11100), .b(g853), .a(g10950) );
  and2_324 AND2_1230 ( .c(g11235), .b(g4529), .a(n1352) );
  and2_323 AND2_1231 ( .c(g5199), .b(g1068), .a(n1161) );
  and2_322 AND2_1232 ( .c(g6316), .b(g1270), .a(n1322) );
  and2_321 AND2_1233 ( .c(g7515), .b(n1384), .a(g70) );
  and2_320 AND2_1234 ( .c(g10583), .b(g10518), .a(g10515) );
  and2_319 AND2_1235 ( .c(g5781), .b(g1537), .a(n1229) );
  and2_318 AND2_1236 ( .c(g8018), .b(g7742), .a(n1245) );
  and2_317 AND2_1237 ( .c(g4401), .b(g1845), .a(g3772) );
  and3_5 AND3_44 ( .d(g8994), .c(n1283), .b(n1307), .a(n1255) );
  and2_316 AND2_1238 ( .c(g2950), .b(n1103), .a(g1666) );
  and2_315 AND2_1239 ( .c(g5510), .b(g1630), .a(n1380) );
  and2_314 AND2_1240 ( .c(g6347), .b(g275), .a(n1221) );
  and2_313 AND2_1241 ( .c(g9357), .b(g962), .a(n1324) );
  and2_312 AND2_1242 ( .c(g4828), .b(g4106), .a(g695) );
  and2_311 AND2_1243 ( .c(g11407), .b(g11249), .a(n1322) );
  and2_310 AND2_1244 ( .c(g4727), .b(g386), .a(g109) );
  and2_309 AND2_1245 ( .c(g10357), .b(n1219), .a(g109) );
  and2_308 AND2_1246 ( .c(g10743), .b(g10639), .a(n1363) );
  and2_307 AND2_1247 ( .c(g5259), .b(g627), .a(n1263) );
  and2_306 AND2_1248 ( .c(g5694), .b(g162), .a(g5361) );
  and2_305 AND2_1249 ( .c(g10769), .b(g10652), .a(n1363) );
  and2_304 AND2_1250 ( .c(g11584), .b(g1318), .a(n1198) );
  and2_303 AND2_1251 ( .c(g4932), .b(g1065), .a(n1380) );
  and2_302 AND2_1252 ( .c(g10768), .b(g10649), .a(n1363) );
  and2_301 AND2_1253 ( .c(g6820), .b(g1362), .a(g5354) );
  and2_300 AND2_1254 ( .c(g4068), .b(g1801), .a(g2276) );
  and2_299 AND2_1255 ( .c(g6317), .b(g1304), .a(n1322) );
  and2_298 AND2_1256 ( .c(g5215), .b(g4276), .a(g3400) );
  and2_297 AND2_1257 ( .c(g4576), .b(g530), .a(g109) );
  and2_296 AND2_1258 ( .c(g4866), .b(g231), .a(g2355) );
  and2_295 AND2_1259 ( .c(g6775), .b(g822), .a(g6231) );
  and2_294 AND2_1260 ( .c(g3829), .b(n1132), .a(g1696) );
  and2_293 AND2_1261 ( .c(g10662), .b(n1224), .a(g10396) );
  and2_292 AND2_1262 ( .c(g8101), .b(g5484), .a(g6740) );
  and2_291 AND2_1263 ( .c(g5825), .b(g3204), .a(g5318) );
  and4_2 AND4_14 ( .e(I6310), .d(n1060), .c(n1143), .b(n1153), .a(n1139) );
  and2_290 AND2_1264 ( .c(g7884), .b(g7457), .a(n1253) );
  and2_289 AND2_1265 ( .c(g5008), .b(g1292), .a(g109) );
  and2_288 AND2_1266 ( .c(g3974), .b(g231), .a(g2355) );
  and2_287 AND2_1267 ( .c(g9949), .b(g9929), .a(n1321) );
  and2_286 AND2_1268 ( .c(g2531), .b(g658), .a(g668) );
  and2_285 AND2_1269 ( .c(g9292), .b(g8878), .a(g48) );
  and2_284 AND2_1270 ( .c(g10778), .b(g1027), .a(g10522) );
  and2_283 AND2_1271 ( .c(g8041), .b(g7524), .a(g5128) );
  and2_282 AND2_1272 ( .c(g6079), .b(g1053), .a(g85) );
  and2_281 AND2_1273 ( .c(g7235), .b(g6663), .a(n1276) );
  and2_280 AND2_1274 ( .c(g9603), .b(g1173), .a(g9125) );
  and2_279 AND2_1275 ( .c(g6840), .b(g248), .a(g5354) );
  and2_278 AND2_1276 ( .c(g9850), .b(g9726), .a(g9560) );
  and2_277 AND2_1277 ( .c(g7988), .b(g1878), .a(g6740) );
  and2_276 AND2_1278 ( .c(g5228), .b(g1086), .a(n1161) );
  and2_275 AND2_1279 ( .c(g7134), .b(g5587), .a(n1236) );
  and2_274 AND2_1280 ( .c(g5934), .b(g5215), .a(n1134) );
  and2_273 AND2_1281 ( .c(g5230), .b(g1265), .a(g109) );
  and2_272 AND2_1282 ( .c(g8168), .b(g34), .a(n1173) );
  and2_271 AND2_1283 ( .c(g9583), .b(g886), .a(g8995) );
  and2_270 AND2_1284 ( .c(g10672), .b(g10414), .a(n1224) );
  and2_269 AND2_1285 ( .c(g3287), .b(g802), .a(g2534) );
  and2_268 AND2_1286 ( .c(g8772), .b(g8627), .a(g5151) );
  and2_267 AND2_1287 ( .c(g4893), .b(g635), .a(n1263) );
  and2_266 AND2_1288 ( .c(g10331), .b(n1214), .a(g109) );
  and2_265 AND2_1289 ( .c(g8505), .b(g8309), .a(g2355) );
  and2_264 AND2_1290 ( .c(g10449), .b(g10420), .a(n1071) );
  and2_263 AND2_1291 ( .c(g11273), .b(g4765), .a(n1357) );
  and2_262 AND2_1292 ( .c(g8734), .b(g8187), .a(n1384) );
  and2_261 AND2_1293 ( .c(g5913), .b(g1041), .a(g85) );
  and2_260 AND2_1294 ( .c(g10448), .b(n1203), .a(n1071) );
  and2_259 AND2_1295 ( .c(g6163), .b(g4572), .a(g5354) );
  and2_258 AND2_1296 ( .c(g6363), .b(g284), .a(n1221) );
  and2_257 AND2_1297 ( .c(g7202), .b(g5226), .a(n1277) );
  and2_256 AND2_1298 ( .c(g11463), .b(g11229), .a(g4421) );
  and2_255 AND2_1299 ( .c(g8074), .b(g718), .a(n1251) );
  and2_254 AND2_1300 ( .c(g4325), .b(g1166), .a(g109) );
  and2_253 AND2_1301 ( .c(g8474), .b(g8383), .a(g3041) );
  and2_252 AND2_1302 ( .c(g11234), .b(g4518), .a(n1353) );
  and2_251 AND2_1303 ( .c(g5266), .b(g718), .a(g3041) );
  and2_250 AND2_1304 ( .c(g4483), .b(g336), .a(g3586) );
  and2_249 AND2_1305 ( .c(g5248), .b(g673), .a(g3041) );
  and2_248 AND2_1306 ( .c(g11514), .b(g11491), .a(g5151) );
  and2_247 AND2_1307 ( .c(g5255), .b(g682), .a(g3041) );
  and2_246 AND2_1308 ( .c(g4106), .b(g3284), .a(g686) );
  and2_245 AND2_1309 ( .c(g2760), .b(g981), .a(g2091) );
  and2_244 AND2_1310 ( .c(g5097), .b(g1786), .a(n1202) );
  and2_243 AND2_1311 ( .c(g5726), .b(g1601), .a(n1215) );
  and2_242 AND2_1312 ( .c(g5497), .b(g560), .a(n1390) );
  and2_241 AND2_1313 ( .c(g5354), .b(g109), .a(n1295) );
  and2_240 AND2_1314 ( .c(g7933), .b(g55), .a(n1383) );
  and2_239 AND2_1315 ( .c(g9617), .b(g9), .a(n1323) );
  and2_238 AND2_1316 ( .c(g9906), .b(g9873), .a(g9683) );
  and2_237 AND2_1317 ( .c(g11012), .b(g5196), .a(n1349) );
  and2_236 AND2_1318 ( .c(g7050), .b(g5001), .a(n1199) );
  and2_235 AND2_1319 ( .c(g10971), .b(g10849), .a(n1142) );
  and2_234 AND2_1320 ( .c(g4904), .b(g1850), .a(n1288) );
  and2_233 AND2_1321 ( .c(g10369), .b(n1187), .a(n1071) );
  and2_232 AND2_1322 ( .c(g8400), .b(g5271), .a(g7101) );
  and2_231 AND2_1323 ( .c(g4345), .b(g1169), .a(n1380) );
  and2_230 AND2_1324 ( .c(g2161), .b(I5084), .a(I5085) );
  and2_229 AND2_1325 ( .c(g5001), .b(g1300), .a(g109) );
  and2_228 AND2_1326 ( .c(g9945), .b(g9925), .a(n1321) );
  and2_227 AND2_1327 ( .c(g7271), .b(g5028), .a(n1236) );
  and2_226 AND2_1328 ( .c(g9709), .b(g1524), .a(n1207) );
  and2_225 AND2_1329 ( .c(g4223), .b(g1003), .a(n1381) );
  and2_224 AND2_1330 ( .c(g10716), .b(g10497), .a(g10396) );
  and2_223 AND2_1331 ( .c(g11291), .b(g11247), .a(n1208) );
  and2_222 AND2_1332 ( .c(g6661), .b(g73), .a(n1176) );
  and2_221 AND2_1333 ( .c(g11173), .b(g491), .a(n1349) );
  and2_220 AND2_1334 ( .c(g6075), .b(g549), .a(n1381) );
  and2_219 AND2_1335 ( .c(g8023), .b(g7367), .a(n1245) );
  and2_218 AND2_1336 ( .c(g9907), .b(g9888), .a(g9686) );
  and2_217 AND2_1337 ( .c(g10582), .b(g10339), .a(n1224) );
  and2_216 AND2_1338 ( .c(g5746), .b(g1589), .a(n1215) );
  and2_215 AND2_1339 ( .c(g5221), .b(g1260), .a(g109) );
  and2_214 AND2_1340 ( .c(g9959), .b(g9950), .a(n1319) );
  and2_213 AND2_1341 ( .c(g7674), .b(g5857), .a(g3880) );
  and2_212 AND2_1342 ( .c(g9690), .b(g266), .a(n1171) );
  and2_211 AND2_1343 ( .c(g6627), .b(g58), .a(n1176) );
  and2_210 AND2_1344 ( .c(g5703), .b(g174), .a(g5361) );
  and2_209 AND2_1345 ( .c(g4522), .b(g360), .a(g3586) );
  and2_208 AND2_1346 ( .c(g4115), .b(g1776), .a(n1103) );
  and2_207 AND2_1347 ( .c(g7541), .b(g7075), .a(n1083) );
  and2_206 AND2_1348 ( .c(g10627), .b(g10452), .a(n1159) );
  and2_205 AND2_1349 ( .c(g4047), .b(n1339), .a(g2276) );
  and2_204 AND2_1350 ( .c(g6526), .b(g76), .a(n1176) );
  and2_203 AND2_1351 ( .c(g2944), .b(n1103), .a(g1669) );
  and2_202 AND2_1352 ( .c(g6646), .b(g360), .a(n1176) );
  and2_201 AND2_1353 ( .c(g7132), .b(g5182), .a(n1199) );
  and2_200 AND2_1354 ( .c(g11029), .b(g401), .a(n1349) );
  and2_199 AND2_1355 ( .c(g8051), .b(g7572), .a(g5128) );
  and2_198 AND2_1356 ( .c(g8127), .b(g1927), .a(n1210) );
  and2_197 AND2_1357 ( .c(g7209), .b(g3804), .a(n1276) );
  and2_196 AND2_1358 ( .c(g11028), .b(g396), .a(n1349) );
  and2_195 AND2_1359 ( .c(g6439), .b(g3631), .a(g5919) );
  and2_194 AND2_1360 ( .c(g10742), .b(g10655), .a(g3586) );
  and2_193 AND2_1361 ( .c(g9110), .b(g8880), .a(g2355) );
  and2_192 AND2_1362 ( .c(g10681), .b(g10567), .a(g3586) );
  and2_191 AND2_1363 ( .c(g4537), .b(g444), .a(g109) );
  and2_190 AND2_1364 ( .c(g9663), .b(g959), .a(n1324) );
  and2_189 AND2_1365 ( .c(g5349), .b(n1158), .a(g4617) );
  and2_188 AND2_1366 ( .c(g8732), .b(g8200), .a(n1384) );
  and2_187 AND2_1367 ( .c(g3807), .b(g3003), .a(g3062) );
  and2_186 AND2_1368 ( .c(g8753), .b(n1231), .a(g8451) );
  and2_185 AND2_1369 ( .c(g5848), .b(g3860), .a(g3661) );
  and2_184 AND2_1370 ( .c(g8508), .b(g8411), .a(g7638) );
  and2_183 AND2_1371 ( .c(g8072), .b(g700), .a(n1251) );
  and2_182 AND2_1372 ( .c(g5699), .b(g1592), .a(n1215) );
  and2_181 AND2_1373 ( .c(g11240), .b(g4560), .a(n1353) );
  and2_180 AND2_1374 ( .c(g5398), .b(g4610), .a(n1048) );
  and2_179 AND2_1375 ( .c(g6616), .b(g6105), .a(n1083) );
  and2_178 AND2_1376 ( .c(g10690), .b(n1201), .a(g3863) );
  and2_177 AND2_1377 ( .c(g8043), .b(g7582), .a(g5128) );
  and2_176 AND2_1378 ( .c(g9590), .b(g895), .a(g8995) );
  and2_175 AND2_1379 ( .c(g4128), .b(n1157), .a(g627) );
  and2_174 AND2_1380 ( .c(g6404), .b(g2132), .a(g5013) );
  and2_173 AND2_1381 ( .c(g6647), .b(g87), .a(n1316) );
  and2_172 AND2_1382 ( .c(g10504), .b(g10001), .a(n1337) );
  and2_171 AND2_1383 ( .c(g9657), .b(g919), .a(g9205) );
  and2_170 AND2_1384 ( .c(g4542), .b(g366), .a(g3586) );
  and2_169 AND2_1385 ( .c(g4330), .b(g1163), .a(g109) );
  and2_168 AND2_1386 ( .c(g3497), .b(g2804), .a(g1900) );
  and2_167 AND2_1387 ( .c(g5524), .b(g1678), .a(n1381) );
  and2_166 AND2_1388 ( .c(g8147), .b(g928), .a(n1209) );
  and2_165 AND2_1389 ( .c(g4554), .b(g542), .a(g109) );
  and2_164 AND2_1390 ( .c(g9899), .b(g9713), .a(n1320) );
  and2_163 AND2_1391 ( .c(g5258), .b(g700), .a(g3041) );
  and2_162 AND2_1392 ( .c(g7736), .b(g5814), .a(g3880) );
  and2_161 AND2_1393 ( .c(g6224), .b(g1520), .a(g5151) );
  and2_160 AND2_1394 ( .c(g10626), .b(g10453), .a(n1159) );
  and2_159 AND2_1395 ( .c(g6320), .b(g1292), .a(n1322) );
  and2_158 AND2_1396 ( .c(g7623), .b(g664), .a(g6488) );
  and2_157 AND2_1397 ( .c(g10299), .b(n1224), .a(g10013) );
  and2_156 AND2_1398 ( .c(g7889), .b(g5304), .a(n1390) );
  and2_155 AND2_1399 ( .c(g10298), .b(n1224), .a(g10007) );
  and2_154 AND2_1400 ( .c(g8413), .b(g722), .a(n1211) );
  and2_153 AND2_1401 ( .c(g3979), .b(g237), .a(g2355) );
  and2_152 AND2_1402 ( .c(g4902), .b(g1848), .a(n1288) );
  and2_151 AND2_1403 ( .c(g5211), .b(g1080), .a(n1161) );
  and2_150 AND2_1404 ( .c(g4512), .b(g357), .a(g3586) );
  and2_149 AND2_1405 ( .c(g7722), .b(g7127), .a(n1276) );
  and2_148 AND2_1406 ( .c(g9844), .b(g9714), .a(g9522) );
  and2_147 AND2_1407 ( .c(g4490), .b(g1141), .a(g109) );
  and2_146 AND2_1408 ( .c(g4823), .b(g207), .a(g2355) );
  and2_145 AND2_1409 ( .c(g6516), .b(g5993), .a(n1083) );
  and2_144 AND2_1410 ( .c(g5026), .b(g1453), .a(g4640) );
  and2_143 AND2_1411 ( .c(g8820), .b(g8705), .a(g3041) );
  and2_142 AND2_1412 ( .c(g10737), .b(g10597), .a(n1363) );
  and3_4 AND3_45 ( .d(g8936), .c(n1273), .b(n1307), .a(n1274) );
  and2_141 AND2_1413 ( .c(g10232), .b(n1224), .a(g9974) );
  and2_140 AND2_1414 ( .c(g6771), .b(g263), .a(n1221) );
  and2_139 AND2_1415 ( .c(g5170), .b(g1811), .a(n1202) );
  and2_138 AND2_1416 ( .c(g8117), .b(g5514), .a(g6740) );
  and2_137 AND2_1417 ( .c(g4529), .b(g448), .a(g109) );
  and2_136 AND2_1418 ( .c(g4348), .b(g3497), .a(g1909) );
  and2_135 AND2_1419 ( .c(g9966), .b(g9956), .a(n1319) );
  and2_134 AND2_1420 ( .c(g5280), .b(n1262), .a(n1116) );
  and2_133 AND2_1421 ( .c(g7139), .b(g5212), .a(n1199) );
  and2_132 AND2_1422 ( .c(g11099), .b(g382), .a(n1163) );
  and2_131 AND2_1423 ( .c(g6892), .b(g6472), .a(g5013) );
  and2_130 AND2_1424 ( .c(g9705), .b(g1580), .a(n1190) );
  and2_129 AND2_1425 ( .c(g10512), .b(g10025), .a(n1337) );
  and2_128 AND2_1426 ( .c(g11098), .b(g849), .a(g10950) );
  and2_127 AND2_1427 ( .c(g8775), .b(g8628), .a(g5151) );
  and2_126 AND2_1428 ( .c(g5083), .b(g2510), .a(n1227) );
  and2_125 AND2_1429 ( .c(g5544), .b(g1687), .a(n1381) );
  and2_124 AND2_1430 ( .c(g11272), .b(g4760), .a(n1356) );
  and2_123 AND2_1431 ( .c(g5483), .b(g1621), .a(n1382) );
  and2_122 AND2_1432 ( .c(g9948), .b(g9928), .a(n1321) );
  and2_121 AND2_1433 ( .c(g4063), .b(g1796), .a(g2276) );
  and2_120 AND2_1434 ( .c(g11462), .b(g11227), .a(g4421) );
  and2_119 AND2_1435 ( .c(g6738), .b(g2531), .a(g5557) );
  and2_118 AND2_1436 ( .c(g8060), .b(g7593), .a(g5919) );
  and2_117 AND2_1437 ( .c(g6244), .b(g1411), .a(g5151) );
  and2_116 AND2_1438 ( .c(g11032), .b(g416), .a(n1349) );
  and2_115 AND2_1439 ( .c(g10445), .b(g9974), .a(n1337) );
  and2_114 AND2_1440 ( .c(g9150), .b(g8882), .a(g2355) );
  and2_113 AND2_1441 ( .c(g10316), .b(g10025), .a(g8574) );
  and2_112 AND2_1442 ( .c(g5756), .b(g1531), .a(n1229) );
  and2_111 AND2_1443 ( .c(g4720), .b(g1023), .a(n1382) );
  and2_110 AND2_1444 ( .c(g9409), .b(g1721), .a(g9052) );
  and2_109 AND2_1445 ( .c(g8995), .b(g48), .a(g8929) );
  and2_108 AND2_1446 ( .c(g6876), .b(g4070), .a(n1267) );
  and2_107 AND2_1447 ( .c(g4989), .b(g1424), .a(g4682) );
  and2_106 AND2_1448 ( .c(g9836), .b(g9737), .a(g9785) );
  and3_3 AND3_46 ( .d(g6656), .c(g109), .b(g6061), .a(n1295) );
  and2_105 AND2_1449 ( .c(g5514), .b(g1941), .a(g3209) );
  and2_104 AND2_1450 ( .c(g8390), .b(g8268), .a(g6465) );
  and2_103 AND2_1451 ( .c(g5003), .b(g1466), .a(g4640) );
  and2_102 AND2_1452 ( .c(g9967), .b(g9957), .a(n1319) );
  and2_101 AND2_1453 ( .c(g5145), .b(g1639), .a(n1382) );
  and2_100 AND2_1454 ( .c(g4834), .b(g219), .a(g2355) );
  and2_99 AND2_1455 ( .c(g4971), .b(g1419), .a(g4682) );
  and2_98 AND2_1456 ( .c(g10753), .b(g10649), .a(n1363) );
  and2_97 AND2_1457 ( .c(g5695), .b(g166), .a(g5361) );
  and2_96 AND2_1458 ( .c(g7613), .b(g6940), .a(g5013) );
  and2_95 AND2_1459 ( .c(g10736), .b(g10658), .a(n1363) );
  and2_94 AND2_1460 ( .c(g11220), .b(g962), .a(n1177) );
  and2_93 AND2_1461 ( .c(g7444), .b(g7277), .a(g5557) );
  and2_92 AND2_1462 ( .c(g5536), .b(g2970), .a(n1286) );
  and2_91 AND2_1463 ( .c(g6663), .b(g6064), .a(n1047) );
  and2_90 AND2_1464 ( .c(g4670), .b(g192), .a(g2355) );
  and2_89 AND2_1465 ( .c(g6824), .b(g1371), .a(g5354) );
  and2_88 AND2_1466 ( .c(g4253), .b(g1074), .a(n1363) );
  and2_87 AND2_1467 ( .c(g8250), .b(g932), .a(n1209) );
  and2_86 AND2_1468 ( .c(g8163), .b(g7960), .a(g636) );
  and2_85 AND2_1469 ( .c(g10764), .b(g10643), .a(n1363) );
  and2_84 AND2_1470 ( .c(g5757), .b(g1552), .a(n1229) );
  and2_83 AND2_1471 ( .c(g10365), .b(g9995), .a(n1337) );
  and2_82 AND2_1472 ( .c(g8032), .b(g7385), .a(n1245) );
  and2_81 AND2_1473 ( .c(g11591), .b(g2988), .a(g11561) );
  and2_80 AND2_1474 ( .c(g8053), .b(g7583), .a(g5919) );
  and2_79 AND2_1475 ( .c(g11147), .b(g321), .a(n1356) );
  and2_78 AND2_1476 ( .c(g5522), .b(g1633), .a(n1382) );
  and2_77 AND2_1477 ( .c(g5115), .b(g1394), .a(g4572) );
  and2_76 AND2_1478 ( .c(g9837), .b(g9697), .a(g9751) );
  and2_75 AND2_1479 ( .c(g9620), .b(g976), .a(n1330) );
  and2_74 AND2_1480 ( .c(g11151), .b(g327), .a(n1356) );
  and2_73 AND2_1481 ( .c(g11172), .b(g486), .a(n1349) );
  and2_72 AND2_1482 ( .c(g7885), .b(g5300), .a(n1391) );
  and2_71 AND2_1483 ( .c(g6064), .b(g5398), .a(n1058) );
  and3_2 AND3_47 ( .d(g8929), .c(n1258), .b(n1307), .a(n1266) );
  and2_70 AND2_1484 ( .c(g5595), .b(g1621), .a(n1388) );
  and2_69 AND2_1485 ( .c(g5537), .b(g2260), .a(n1277) );
  and2_68 AND2_1486 ( .c(g9842), .b(g9708), .a(g9516) );
  and2_67 AND2_1487 ( .c(g4141), .b(g1791), .a(n1103) );
  and2_66 AND2_1488 ( .c(g4341), .b(g339), .a(g3586) );
  and2_65 AND2_1489 ( .c(g9192), .b(g48), .a(g8955) );
  and2_64 AND2_1490 ( .c(g7679), .b(g1950), .a(n1257) );
  and2_63 AND2_1491 ( .c(g7378), .b(g5847), .a(g3880) );
  and2_62 AND2_1492 ( .c(g5612), .b(g1627), .a(n1390) );
  and2_61 AND2_1493 ( .c(g3939), .b(g213), .a(g2355) );
  and2_60 AND2_1494 ( .c(g7135), .b(g869), .a(g6355) );
  and2_59 AND2_1495 ( .c(g10970), .b(n1193), .a(g1811) );
  and2_58 AND2_1496 ( .c(g11025), .b(g426), .a(n1349) );
  and2_57 AND2_1497 ( .c(g9854), .b(g9730), .a(g9566) );
  and2_56 AND2_1498 ( .c(g7182), .b(g1878), .a(g6003) );
  and2_55 AND2_1499 ( .c(g9941), .b(g9921), .a(n1320) );
  and2_54 AND2_1500 ( .c(g6194), .b(g554), .a(n1382) );
  and2_53 AND2_1501 ( .c(g5128), .b(n1295), .a(g109) );
  and2_52 AND2_1502 ( .c(g4962), .b(g1651), .a(n1202) );
  and2_51 AND2_1503 ( .c(g4358), .b(g1209), .a(n1382) );
  and2_50 AND2_1504 ( .c(g8683), .b(g4803), .a(g8549) );
  and2_49 AND2_1505 ( .c(g4506), .b(g1113), .a(g109) );
  and2_48 AND2_1506 ( .c(g6471), .b(g5224), .a(n1216) );
  and2_47 AND2_1507 ( .c(g8778), .b(n1261), .a(n1055) );
  and2_46 AND2_1508 ( .c(g11281), .b(g4788), .a(n1356) );
  and2_45 AND2_1509 ( .c(g8735), .b(n1231), .a(g8451) );
  and2_44 AND2_1510 ( .c(g11146), .b(g318), .a(n1357) );
  and2_43 AND2_1511 ( .c(g3904), .b(g2948), .a(g627) );
  and2_42 AND2_1512 ( .c(g8075), .b(g727), .a(n1251) );
  and2_41 AND2_1513 ( .c(g9829), .b(g9723), .a(g9785) );
  and3_1 AND3_48 ( .d(g8949), .c(n1259), .b(n1307), .a(n1266) );
  and2_40 AND2_1514 ( .c(g7632), .b(g7184), .a(n1240) );
  and2_39 AND2_1515 ( .c(g11290), .b(g11246), .a(n1208) );
  and2_38 AND2_1516 ( .c(g6350), .b(g5837), .a(n1363) );
  and2_37 AND2_1517 ( .c(g10599), .b(g10448), .a(n1159) );
  and2_36 AND2_1518 ( .c(g5902), .b(g2555), .a(g4977) );
  and4_1 AND4_15 ( .e(I6337), .d(g201), .c(n1153), .b(n1143), .a(n1060) );
  and2_35 AND2_1519 ( .c(g2276), .b(g1765), .a(g1610) );
  and2_34 AND2_1520 ( .c(g6438), .b(g5853), .a(g5013) );
  and2_33 AND2_1521 ( .c(g5512), .b(g1660), .a(n1161) );
  and2_32 AND2_1522 ( .c(g5090), .b(n1339), .a(n1202) );
  and2_31 AND2_1523 ( .c(g7719), .b(g718), .a(g6488) );
  and2_30 AND2_1524 ( .c(g2561), .b(g742), .a(g741) );
  and2_29 AND2_1525 ( .c(g3695), .b(g1712), .a(n1363) );
  and2_28 AND2_1526 ( .c(g8603), .b(n1278), .a(n1205) );
  and2_27 AND2_1527 ( .c(g8039), .b(g7587), .a(g5128) );
  and2_26 AND2_1528 ( .c(g9610), .b(g925), .a(g9192) );
  and2_25 AND2_1529 ( .c(g3536), .b(g1289), .a(n1110) );
  and2_24 AND2_1530 ( .c(g5529), .b(g2257), .a(n1286) );
  and2_23 AND2_1531 ( .c(g5148), .b(g1107), .a(n1235) );
  and2_22 AND2_1532 ( .c(g9124), .b(g8881), .a(g2355) );
  and2_21 AND2_1533 ( .c(g9324), .b(g8879), .a(g48) );
  and2_20 AND2_1534 ( .c(g4559), .b(n1067), .a(g3829) );
  and2_19 AND2_1535 ( .c(g10561), .b(g10549), .a(n1159) );
  and2_18 AND2_1536 ( .c(g5698), .b(g1571), .a(n1215) );
  and2_17 AND2_1537 ( .c(g11226), .b(n1332), .a(n1191) );
  and2_16 AND2_1538 ( .c(g10295), .b(n1224), .a(g9995) );
  and2_15 AND2_1539 ( .c(g5260), .b(g1092), .a(n1161) );
  and2_14 AND2_1540 ( .c(g10680), .b(g10564), .a(g3586) );
  and2_13 AND2_1541 ( .c(g6822), .b(g231), .a(g5354) );
  and2_12 AND2_1542 ( .c(g4905), .b(g1853), .a(n1288) );
  and2_11 AND2_1543 ( .c(g11551), .b(g11538), .a(n1365) );
  and2_10 AND2_1544 ( .c(g3047), .b(g1227), .a(g2306) );
  and2_9 AND2_1545 ( .c(g9849), .b(g293), .a(g9313) );
  and2_8 AND2_1546 ( .c(g5279), .b(n1333), .a(n1202) );
  and2_7 AND2_1547 ( .c(g8404), .b(g686), .a(n1211) );
  and2_6 AND2_1548 ( .c(g5720), .b(g170), .a(g5361) );
  and2_5 AND2_1549 ( .c(g5318), .b(g4401), .a(g1857) );
  and2_4 AND2_1550 ( .c(g8764), .b(n1231), .a(g8451) );
  and2_3 AND2_1551 ( .c(g11376), .b(g11318), .a(n1223) );
  and2_2 AND2_1552 ( .c(g11297), .b(g4565), .a(n1357) );
  and2_1 AND2_1553 ( .c(g9898), .b(g9710), .a(n1320) );
  or2_0 OR2_0 ( .c(g6895), .b(g6776), .a(g4875) );
  or2_586 OR2_1 ( .c(g7189), .b(g6632), .a(g4421) );
  or2_585 OR2_2 ( .c(g9510), .b(g9125), .a(g9111) );
  or2_584 OR2_3 ( .c(g7297), .b(g7132), .a(g6323) );
  or2_583 OR2_4 ( .c(g9088), .b(g8927), .a(g41) );
  or2_582 OR2_5 ( .c(g9923), .b(g9865), .a(g9707) );
  or2_581 OR2_6 ( .c(g6485), .b(g5848), .a(g5067) );
  or2_580 OR2_7 ( .c(g8771), .b(g5483), .a(g8652) );
  or2_579 OR2_8 ( .c(g5813), .b(g5617), .a(g4869) );
  or2_578 OR2_9 ( .c(g7963), .b(n1253), .a(g7182) );
  or2_577 OR2_10 ( .c(g10643), .b(g10624), .a(g7736) );
  or3_0 OR3_0 ( .d(g9886), .c(g9607), .b(g9592), .a(g9759) );
  or3_61 OR3_1 ( .d(g9951), .c(g9902), .b(g9899), .a(g9803) );
  or2_576 OR2_11 ( .c(g11625), .b(g6535), .a(g11597) );
  or2_575 OR2_12 ( .c(g8945), .b(g8801), .a(g8710) );
  or2_574 OR2_13 ( .c(g10489), .b(g1718), .a(g10367) );
  or2_573 OR2_14 ( .c(g10559), .b(g4141), .a(g10512) );
  or2_572 OR2_15 ( .c(g10558), .b(g4126), .a(g10510) );
  or2_571 OR2_16 ( .c(g11338), .b(g11283), .a(g11178) );
  or2_570 OR2_17 ( .c(g8435), .b(g8403), .a(g8075) );
  or2_569 OR2_18 ( .c(g10544), .b(g1718), .a(g10495) );
  or2_568 OR2_19 ( .c(g6911), .b(g6342), .a(g5681) );
  or2_567 OR2_20 ( .c(g10865), .b(g5538), .a(g10752) );
  or2_566 OR2_21 ( .c(g3698), .b(n1392), .a(g869) );
  or2_565 OR2_22 ( .c(g8214), .b(g7472), .a(g82) );
  or2_564 OR2_23 ( .c(g6124), .b(g5181), .a(g5188) );
  or2_563 OR2_24 ( .c(g6469), .b(g5698), .a(g4959) );
  or2_562 OR2_25 ( .c(g5587), .b(g4714), .a(g3904) );
  or2_561 OR2_26 ( .c(g6177), .b(g5444), .a(g4712) );
  or3_60 OR3_2 ( .d(I14585), .c(g8995), .b(g9205), .a(g9192) );
  or2_560 OR2_27 ( .c(g9891), .b(n1327), .a(n1182) );
  or2_559 OR2_28 ( .c(g9913), .b(g9849), .a(g9691) );
  or4_0 OR4_0 ( .e(I5600), .d(g496), .c(g491), .b(g486), .a(g481) );
  or2_558 OR2_29 ( .c(g11257), .b(g11234), .a(g11019) );
  or2_557 OR2_30 ( .c(g8236), .b(g7526), .a(g82) );
  or2_556 OR2_31 ( .c(g7385), .b(g7235), .a(g6746) );
  or2_555 OR2_32 ( .c(g6898), .b(g6790), .a(g4881) );
  or2_554 OR2_33 ( .c(g6900), .b(g6787), .a(g6246) );
  or2_553 OR2_34 ( .c(g4264), .b(g4048), .a(g4053) );
  or3_59 OR3_3 ( .d(g9726), .c(g9411), .b(g9420), .a(g9489) );
  or2_552 OR2_35 ( .c(g6088), .b(g5260), .a(g4522) );
  or2_551 OR2_36 ( .c(g6923), .b(g6353), .a(g5695) );
  or2_550 OR2_37 ( .c(g8194), .b(g5168), .a(g7940) );
  or3_58 OR3_4 ( .d(g9676), .c(n1327), .b(n1331), .a(n1323) );
  or2_549 OR2_38 ( .c(g11256), .b(g11186), .a(g11018) );
  or2_548 OR2_39 ( .c(g3860), .b(g3107), .a(g2167) );
  or2_547 OR2_40 ( .c(g11280), .b(g11254), .a(g11153) );
  or4_60 OR4_1 ( .e(g9727), .d(g9650), .c(g9663), .b(g9362), .a(I14866) );
  or2_546 OR2_41 ( .c(g4997), .b(g4581), .a(g4584) );
  or2_545 OR2_42 ( .c(g11624), .b(g11595), .a(g11571) );
  or2_544 OR2_43 ( .c(g11300), .b(g11213), .a(g11091) );
  or2_543 OR2_44 ( .c(g4238), .b(g3999), .a(g4007) );
  or2_542 OR2_45 ( .c(g8814), .b(g7945), .a(g8728) );
  or2_541 OR2_46 ( .c(g10401), .b(g9317), .a(g10291) );
  or2_540 OR2_47 ( .c(g8773), .b(g5491), .a(g8653) );
  or2_539 OR2_48 ( .c(g11231), .b(g11156), .a(g11013) );
  or2_538 OR2_49 ( .c(g10864), .b(g5532), .a(g10751) );
  or2_537 OR2_50 ( .c(g9624), .b(g9316), .a(g9313) );
  or3_57 OR3_5 ( .d(g9953), .c(g9945), .b(g9939), .a(g9669) );
  or2_536 OR2_51 ( .c(g6122), .b(g5172), .a(g5180) );
  or2_535 OR2_52 ( .c(g6465), .b(g5825), .a(g5041) );
  or2_534 OR2_53 ( .c(g6934), .b(g6363), .a(g5720) );
  or2_533 OR2_54 ( .c(g7664), .b(g6855), .a(n1392) );
  or2_532 OR2_55 ( .c(g7246), .b(g6465), .a(g6003) );
  or2_531 OR2_56 ( .c(g7203), .b(g6640), .a(g6058) );
  or2_530 OR2_57 ( .c(g6096), .b(g5268), .a(g4542) );
  or2_529 OR2_58 ( .c(g9747), .b(n1328), .a(g9509) );
  or2_528 OR2_59 ( .c(g11314), .b(g11224), .a(g11102) );
  or2_527 OR2_60 ( .c(g10733), .b(g5227), .a(g10522) );
  or2_526 OR2_61 ( .c(g8921), .b(g8827), .a(g8748) );
  or4_59 OR4_2 ( .e(I15054), .d(n1173), .c(n1327), .b(g9624), .a(g9785) );
  or2_525 OR2_62 ( .c(g11269), .b(g11196), .a(g11031) );
  or2_524 OR2_63 ( .c(g5555), .b(g4389), .a(g4397) );
  or2_523 OR2_64 ( .c(g11268), .b(g11194), .a(g11030) );
  or2_522 OR2_65 ( .c(g10485), .b(g9317), .a(g10376) );
  or2_521 OR2_66 ( .c(g10555), .b(g4103), .a(g10504) );
  or2_520 OR2_67 ( .c(g6481), .b(g5722), .a(g4972) );
  or2_519 OR2_68 ( .c(g10712), .b(g10662), .a(g8574) );
  or2_518 OR2_69 ( .c(g11335), .b(g11279), .a(g11175) );
  or2_517 OR2_70 ( .c(g8249), .b(g8018), .a(g7710) );
  or2_516 OR2_71 ( .c(g7638), .b(g7265), .a(g6488) );
  or2_515 OR2_72 ( .c(g10567), .b(g10514), .a(g7378) );
  or2_514 OR2_73 ( .c(g11487), .b(g6662), .a(g11464) );
  or4_58 OR4_3 ( .e(I15210), .d(g9839), .c(g9964), .b(g9852), .a(g9882) );
  or4_57 OR4_4 ( .e(I5805), .d(g2102), .c(g2099), .b(g2096), .a(g2088) );
  or2_513 OR2_74 ( .c(g8941), .b(g8796), .a(g8706) );
  or2_512 OR2_75 ( .c(g11443), .b(g7130), .a(g11407) );
  or2_511 OR2_76 ( .c(g4231), .b(g3991), .a(g3998) );
  or2_510 OR2_77 ( .c(g11278), .b(g11253), .a(g11150) );
  or4_56 OR4_5 ( .e(I15039), .d(n1173), .c(n1327), .b(g9624), .a(g9785) );
  or2_509 OR2_78 ( .c(g11286), .b(g10670), .a(g11209) );
  or2_508 OR2_79 ( .c(g8431), .b(g8387), .a(g8071) );
  or2_507 OR2_80 ( .c(g7133), .b(g6616), .a(g1713) );
  or2_506 OR2_81 ( .c(g11306), .b(g11216), .a(g11095) );
  or2_505 OR2_82 ( .c(g8252), .b(g7988), .a(g7679) );
  or2_504 OR2_83 ( .c(g8812), .b(g7939), .a(g8724) );
  or2_503 OR2_84 ( .c(g7846), .b(g7722), .a(g7241) );
  or2_502 OR2_85 ( .c(g3875), .b(g3275), .a(g12) );
  or2_501 OR2_86 ( .c(g5996), .b(g5473), .a(g3908) );
  or2_500 OR2_87 ( .c(g6592), .b(g5100), .a(g5882) );
  or2_499 OR2_88 ( .c(g8286), .b(g8107), .a(g7823) );
  or2_498 OR2_89 ( .c(g10501), .b(g4161), .a(g10445) );
  or2_497 OR2_90 ( .c(g10728), .b(g4973), .a(g10642) );
  or2_496 OR2_91 ( .c(g8270), .b(g7894), .a(g3434) );
  or2_495 OR2_92 ( .c(g7290), .b(g7046), .a(g6316) );
  or2_494 OR2_93 ( .c(g6068), .b(g5220), .a(g4497) );
  or2_493 OR2_94 ( .c(g6468), .b(g5690), .a(g4950) );
  or2_492 OR2_95 ( .c(g11217), .b(g11144), .a(g11005) );
  or2_491 OR2_96 ( .c(g11478), .b(g6532), .a(g11455) );
  or4_55 OR4_6 ( .e(g9536), .d(g9335), .c(g9331), .b(g9328), .a(g9324) );
  or2_490 OR2_97 ( .c(g5981), .b(g5074), .a(g4383) );
  or2_489 OR2_98 ( .c(g11486), .b(g6654), .a(g11463) );
  or2_488 OR2_99 ( .c(g8377), .b(g8185), .a(g7958) );
  or2_487 OR2_100 ( .c(g8206), .b(g7459), .a(g82) );
  or2_486 OR2_101 ( .c(g11580), .b(g11413), .a(g11544) );
  or2_485 OR2_102 ( .c(g8287), .b(g8117), .a(g7824) );
  or2_484 OR2_103 ( .c(g11223), .b(g11147), .a(g11008) );
  or2_483 OR2_104 ( .c(g9522), .b(n1328), .a(g9125) );
  or2_482 OR2_105 ( .c(g8199), .b(g7902), .a(g7444) );
  or2_481 OR2_106 ( .c(g5802), .b(g5601), .a(g4837) );
  or2_480 OR2_107 ( .c(g11321), .b(g11230), .a(g11105) );
  or2_479 OR2_108 ( .c(g6524), .b(g5746), .a(g4996) );
  or2_478 OR2_109 ( .c(g10664), .b(g10240), .a(g10582) );
  or2_477 OR2_110 ( .c(g7257), .b(g6701), .a(g4725) );
  or2_476 OR2_111 ( .c(g7301), .b(g7140), .a(g6327) );
  or2_475 OR2_112 ( .c(g10484), .b(g9317), .a(n1165) );
  or2_474 OR2_113 ( .c(g10554), .b(g4097), .a(g10503) );
  or2_473 OR2_114 ( .c(g8259), .b(g8028), .a(g7719) );
  or2_472 OR2_115 ( .c(g11334), .b(g11277), .a(g11174) );
  or2_471 OR2_116 ( .c(g8819), .b(g7957), .a(g8734) );
  or2_470 OR2_117 ( .c(g8923), .b(g8846), .a(g8763) );
  or2_469 OR2_118 ( .c(g8488), .b(n1254), .a(g8390) );
  or2_468 OR2_119 ( .c(g7441), .b(g7271), .a(g5867) );
  or2_467 OR2_120 ( .c(g6026), .b(g5507), .a(g3970) );
  or2_466 OR2_121 ( .c(g10799), .b(g6225), .a(g10769) );
  or2_465 OR2_122 ( .c(g10798), .b(g6217), .a(g10768) );
  or2_464 OR2_123 ( .c(g10805), .b(g10759), .a(g10760) );
  or2_463 OR2_124 ( .c(g10732), .b(g4358), .a(g10661) );
  or2_462 OR2_125 ( .c(g6061), .b(g5204), .a(g4) );
  or2_461 OR2_126 ( .c(g9512), .b(n1325), .a(g9125) );
  or2_460 OR2_127 ( .c(g10013), .b(I15214), .a(I15215) );
  or2_459 OR2_128 ( .c(g8806), .b(g7931), .a(g8718) );
  or2_458 OR2_129 ( .c(g8943), .b(g8837), .a(g8749) );
  or2_457 OR2_130 ( .c(g11293), .b(g11211), .a(g10818) );
  or2_456 OR2_131 ( .c(g11265), .b(g11189), .a(g11027) );
  or2_455 OR2_132 ( .c(g8887), .b(g8842), .a(g8755) );
  or2_454 OR2_133 ( .c(g5838), .b(g5612), .a(g4866) );
  or2_453 OR2_134 ( .c(g6514), .b(g5738), .a(g4992) );
  or2_452 OR2_135 ( .c(g8322), .b(g8136), .a(g6891) );
  or2_451 OR2_136 ( .c(g8230), .b(g7515), .a(g82) );
  or2_450 OR2_137 ( .c(g5809), .b(g5611), .a(g4865) );
  or2_449 OR2_138 ( .c(g8433), .b(g8399), .a(g8073) );
  or2_448 OR2_139 ( .c(g11579), .b(g5123), .a(g11551) );
  or2_447 OR2_140 ( .c(g10771), .b(g5533), .a(g10684) );
  or2_446 OR2_141 ( .c(g11615), .b(g11601), .a(g11592) );
  or2_445 OR2_142 ( .c(g9367), .b(g9335), .a(g9331) );
  or3_56 OR3_6 ( .d(g9872), .c(g9617), .b(g9594), .a(g9750) );
  or2_444 OR2_143 ( .c(g6522), .b(g5744), .a(g4994) );
  or2_443 OR2_144 ( .c(g8266), .b(g7885), .a(g3412) );
  or2_442 OR2_145 ( .c(g10414), .b(g10300), .a(g8574) );
  or2_441 OR2_146 ( .c(g11275), .b(g11248), .a(g11148) );
  or2_440 OR2_147 ( .c(g11430), .b(g11387), .a(g4006) );
  or2_439 OR2_148 ( .c(g8248), .b(g8014), .a(g7707) );
  or3_55 OR3_7 ( .d(g9686), .c(n1327), .b(n1331), .a(n1323) );
  or2_438 OR2_149 ( .c(g8815), .b(g7948), .a(g8730) );
  or2_437 OR2_150 ( .c(g7183), .b(g6623), .a(g4421) );
  or2_436 OR2_151 ( .c(g5983), .b(g5084), .a(g4392) );
  or2_435 OR2_152 ( .c(g8154), .b(g7891), .a(g6879) );
  or2_434 OR2_153 ( .c(g6537), .b(g5781), .a(g5005) );
  or2_433 OR2_154 ( .c(g4309), .b(g4069), .a(g4079) );
  or2_432 OR2_155 ( .c(g10725), .b(g4962), .a(g10634) );
  or2_431 OR2_156 ( .c(g6243), .b(g5537), .a(g4144) );
  or4_54 OR4_7 ( .e(I6351), .d(g2405), .c(g2389), .b(g2380), .a(g2372) );
  or3_54 OR3_8 ( .d(g9519), .c(n1328), .b(n1325), .a(g9125) );
  or2_430 OR2_157 ( .c(g9740), .b(g9418), .a(n1340) );
  or2_429 OR2_158 ( .c(g8267), .b(g7889), .a(g3422) );
  or3_53 OR3_9 ( .d(g10744), .c(g10381), .b(n1296), .a(I16427) );
  or2_428 OR2_159 ( .c(g6542), .b(g5789), .a(g5010) );
  or2_427 OR2_160 ( .c(g7303), .b(g7145), .a(g6329) );
  or2_426 OR2_161 ( .c(g10652), .b(g10627), .a(g7743) );
  or2_425 OR2_162 ( .c(g5036), .b(g4871), .a(g4162) );
  or2_424 OR2_163 ( .c(g7240), .b(g6687), .a(g6095) );
  or2_423 OR2_164 ( .c(g8221), .b(g7496), .a(g82) );
  or2_422 OR2_165 ( .c(g6902), .b(g6794), .a(g4223) );
  or3_52 OR3_10 ( .d(I14776), .c(g8995), .b(g9205), .a(g9192) );
  or2_421 OR2_166 ( .c(g10500), .b(g4157), .a(g10442) );
  or2_420 OR2_167 ( .c(g4052), .b(g2862), .a(g2515) );
  or4_53 OR4_8 ( .e(I14858), .d(g9585), .c(g9595), .b(g9610), .a(g9602) );
  or2_419 OR2_168 ( .c(g6529), .b(g5757), .a(g5000) );
  or2_418 OR2_169 ( .c(g11264), .b(g11188), .a(g11026) );
  or4_52 OR4_9 ( .e(I15209), .d(g8169), .c(g9905), .b(g9934), .a(g9830) );
  or2_417 OR2_170 ( .c(g8241), .b(g7536), .a(g82) );
  or2_416 OR2_171 ( .c(g10795), .b(g6199), .a(g10764) );
  or2_415 OR2_172 ( .c(g11607), .b(g11586), .a(g11557) );
  or2_414 OR2_173 ( .c(g8644), .b(g8123), .a(g8464) );
  or3_51 OR3_11 ( .d(g4682), .c(g3563), .b(n1392), .a(g1570) );
  or2_413 OR2_174 ( .c(g8818), .b(g7955), .a(g8733) );
  or2_412 OR2_175 ( .c(g2984), .b(g2528), .a(g2522) );
  or2_411 OR2_176 ( .c(g9931), .b(g8931), .a(g9900) );
  or2_410 OR2_177 ( .c(g3414), .b(g2911), .a(g2917) );
  or2_409 OR2_178 ( .c(g9515), .b(n1328), .a(n1325) );
  or2_408 OR2_179 ( .c(g10724), .b(g10312), .a(g10672) );
  or2_407 OR2_180 ( .c(g7294), .b(g7068), .a(g6320) );
  or2_406 OR2_181 ( .c(g5189), .b(g4345), .a(n1367) );
  or2_405 OR2_182 ( .c(g8614), .b(g8365), .a(g8510) );
  or2_404 OR2_183 ( .c(g3513), .b(g3118), .a(g2180) );
  or2_403 OR2_184 ( .c(g6909), .b(g6346), .a(g5309) );
  or4_51 OR4_10 ( .e(I5571), .d(g396), .c(g391), .b(g386), .a(g426) );
  or2_402 OR2_185 ( .c(g4283), .b(g4059), .a(g4063) );
  or2_401 OR2_186 ( .c(g8939), .b(g8791), .a(g8701) );
  or2_400 OR2_187 ( .c(g2514), .b(I5599), .a(I5600) );
  or2_399 OR2_188 ( .c(g11327), .b(g11297), .a(g11167) );
  or2_398 OR2_189 ( .c(g8187), .b(g7542), .a(g82) );
  or2_397 OR2_190 ( .c(g11606), .b(g11585), .a(g11556) );
  or2_396 OR2_191 ( .c(g11303), .b(g11214), .a(g11092) );
  or2_395 OR2_192 ( .c(g5309), .b(n1254), .a(g4401) );
  or3_50 OR3_12 ( .d(g9528), .c(n1325), .b(g9125), .a(g9111) );
  or2_394 OR2_193 ( .c(g8200), .b(g7535), .a(g82) );
  or3_49 OR3_13 ( .d(g2522), .c(g833), .b(g829), .a(I5629) );
  or4_50 OR4_11 ( .e(g2315), .d(g1163), .c(g1166), .b(g1113), .a(I5363) );
  or2_393 OR2_194 ( .c(g6506), .b(g5731), .a(g4989) );
  or2_392 OR2_195 ( .c(g10649), .b(g10626), .a(g7741) );
  or2_391 OR2_196 ( .c(g8159), .b(g7895), .a(g6886) );
  or2_390 OR2_197 ( .c(g7626), .b(g7060), .a(n1264) );
  or2_389 OR2_198 ( .c(g10770), .b(g5525), .a(g10682) );
  or2_388 OR2_199 ( .c(g9566), .b(g9052), .a(n1329) );
  or2_387 OR2_200 ( .c(g11483), .b(g6633), .a(g11460) );
  or2_386 OR2_201 ( .c(g8811), .b(g7935), .a(g8722) );
  or3_48 OR3_14 ( .d(g8642), .c(g30), .b(g31), .a(n1184) );
  or2_385 OR2_202 ( .c(g6545), .b(g5795), .a(g5025) );
  or2_384 OR2_203 ( .c(g10767), .b(g5500), .a(g10681) );
  or2_383 OR2_204 ( .c(g11326), .b(g11296), .a(g11166) );
  or2_382 OR2_205 ( .c(g10898), .b(g4220), .a(g10777) );
  or2_381 OR2_206 ( .c(g11252), .b(g11099), .a(g10969) );
  or2_380 OR2_207 ( .c(g10719), .b(g10303), .a(g10666) );
  or2_379 OR2_208 ( .c(g4609), .b(g3400), .a(g119) );
  or2_378 OR2_209 ( .c(g6507), .b(g5732), .a(g4990) );
  or2_377 OR2_210 ( .c(g10718), .b(g6238), .a(g10706) );
  or2_376 OR2_211 ( .c(g10521), .b(I16148), .a(I16149) );
  or2_375 OR2_212 ( .c(g7075), .b(g5104), .a(g6530) );
  or2_374 OR2_213 ( .c(g7292), .b(g7055), .a(g6318) );
  or2_373 OR2_214 ( .c(g10861), .b(g5523), .a(g10745) );
  or2_372 OR2_215 ( .c(g8417), .b(g8246), .a(g7721) );
  or2_371 OR2_216 ( .c(g6515), .b(g5739), .a(g4993) );
  or4_49 OR4_12 ( .e(I14855), .d(g9583), .c(g9593), .b(g9601), .a(g9596) );
  or4_48 OR4_13 ( .e(I15205), .d(g9838), .c(g9963), .b(g9850), .a(g9878) );
  or4_47 OR4_14 ( .e(I15051), .d(n1173), .c(g9673), .b(g9624), .a(g9785) );
  or3_47 OR3_15 ( .d(g9724), .c(g9409), .b(g9419), .a(g9615) );
  or2_370 OR2_217 ( .c(g6528), .b(g5756), .a(g4999) );
  or2_369 OR2_218 ( .c(g8823), .b(g8778), .a(g8693) );
  or2_368 OR2_219 ( .c(g7503), .b(g6887), .a(g6430) );
  or2_367 OR2_220 ( .c(g8148), .b(g7884), .a(g6872) );
  or2_366 OR2_221 ( .c(g8649), .b(g8499), .a(n1264) );
  or2_365 OR2_222 ( .c(g3584), .b(g2863), .a(g2516) );
  or2_364 OR2_223 ( .c(g10776), .b(g5544), .a(g10758) );
  or3_46 OR3_16 ( .d(g9680), .c(n1327), .b(n1331), .a(n1323) );
  or2_363 OR2_224 ( .c(g10859), .b(g5512), .a(g10742) );
  or3_45 OR3_17 ( .d(I14866), .c(g9590), .b(g9609), .a(g9619) );
  or2_362 OR2_225 ( .c(g7299), .b(g7138), .a(g6325) );
  or2_361 OR2_226 ( .c(g10858), .b(g5501), .a(g10741) );
  or2_360 OR2_227 ( .c(g8193), .b(g5145), .a(g7937) );
  or3_44 OR3_18 ( .d(g9511), .c(n1325), .b(g9125), .a(g9111) );
  or2_359 OR2_228 ( .c(g7738), .b(g7200), .a(g6738) );
  or2_358 OR2_229 ( .c(g7244), .b(g6699), .a(g4720) );
  or2_357 OR2_230 ( .c(g3425), .b(g2895), .a(g2910) );
  or2_356 OR2_231 ( .c(g7478), .b(g6884), .a(g6423) );
  or3_43 OR3_19 ( .d(g9714), .c(g9664), .b(g9366), .a(g9654) );
  or2_355 OR2_232 ( .c(g10025), .b(I15224), .a(I15225) );
  or2_354 OR2_233 ( .c(g6908), .b(g6345), .a(g4229) );
  or2_353 OR2_234 ( .c(g5028), .b(g4836), .a(g4128) );
  or2_352 OR2_235 ( .c(g8253), .b(g8023), .a(g7718) );
  or2_351 OR2_236 ( .c(g8938), .b(g8789), .a(g8699) );
  or2_350 OR2_237 ( .c(g8813), .b(g7943), .a(g8726) );
  or2_349 OR2_238 ( .c(g9736), .b(g9430), .a(g9416) );
  or2_348 OR2_239 ( .c(g9968), .b(I15171), .a(I15172) );
  or2_347 OR2_240 ( .c(g8552), .b(g8217), .a(g8388) );
  or2_346 OR2_241 ( .c(g5910), .b(g5023), .a(g4341) );
  or2_345 OR2_242 ( .c(g11249), .b(g6162), .a(g11143) );
  or2_344 OR2_243 ( .c(g11482), .b(g6628), .a(g11459) );
  or4_46 OR4_15 ( .e(g9722), .d(g9612), .c(g9643), .b(g9410), .a(I14855) );
  or4_45 OR4_16 ( .e(I15204), .d(g8168), .c(g9904), .b(g9933), .a(g9829) );
  or2_343 OR2_244 ( .c(g7236), .b(g6684), .a(g6092) );
  or3_42 OR3_20 ( .d(I14596), .c(g8995), .b(g9205), .a(g9192) );
  or2_342 OR2_245 ( .c(g8645), .b(g8127), .a(g8469) );
  or2_341 OR2_246 ( .c(g11647), .b(g6622), .a(g11637) );
  or2_340 OR2_247 ( .c(g6777), .b(n1305), .a(g48) );
  or3_41 OR3_21 ( .d(g9737), .c(g9657), .b(g9658), .a(g9655) );
  or4_44 OR4_17 ( .e(I16149), .d(g10472), .c(g10470), .b(g10468), .a(g10467)
         );
  or2_339 OR2_248 ( .c(g11233), .b(g11085), .a(g10946) );
  or2_338 OR2_249 ( .c(g8607), .b(g8406), .a(g8554) );
  or4_43 OR4_18 ( .e(I16148), .d(g10386), .c(g10384), .b(g10476), .a(g10474)
         );
  or2_337 OR2_250 ( .c(g8158), .b(g7893), .a(g6883) );
  or2_336 OR2_251 ( .c(g5846), .b(g4932), .a(g4236) );
  or2_335 OR2_252 ( .c(g5396), .b(g4481), .a(g3684) );
  or2_334 OR2_253 ( .c(g5803), .b(g5575), .a(g4820) );
  or2_333 OR2_254 ( .c(g11331), .b(g11272), .a(g11171) );
  or2_332 OR2_255 ( .c(g7295), .b(g7071), .a(g6321) );
  or2_331 OR2_256 ( .c(g6541), .b(g5788), .a(g5009) );
  or2_330 OR2_257 ( .c(g8615), .b(g8413), .a(g8557) );
  or2_329 OR2_258 ( .c(g9742), .b(n1328), .a(g9528) );
  or2_328 OR2_259 ( .c(g9926), .b(g9868), .a(g9715) );
  or2_327 OR2_260 ( .c(g9754), .b(n1328), .a(g9511) );
  or2_326 OR2_261 ( .c(g8284), .b(g8102), .a(g7821) );
  or2_325 OR2_262 ( .c(g2204), .b(g1393), .a(g1394) );
  or2_324 OR2_263 ( .c(g7471), .b(g6880), .a(g6416) );
  or2_323 OR2_264 ( .c(g7242), .b(g6693), .a(g6098) );
  or2_322 OR2_265 ( .c(g5847), .b(g5626), .a(g4877) );
  or2_321 OR2_266 ( .c(g6901), .b(g6788), .a(g6247) );
  or2_320 OR2_267 ( .c(g8559), .b(g8380), .a(n1254) );
  or3_40 OR3_22 ( .d(g9729), .c(g9618), .b(g9357), .a(g9656) );
  or2_319 OR2_268 ( .c(g10860), .b(g5513), .a(g10743) );
  or2_318 OR2_269 ( .c(g9927), .b(g9869), .a(g9716) );
  or2_317 OR2_270 ( .c(g10497), .b(g48), .a(g10396) );
  or4_42 OR4_19 ( .e(g9885), .d(n1327), .c(g9598), .b(g9662), .a(g9746) );
  or4_41 OR4_20 ( .e(g2528), .d(g861), .c(g857), .b(g853), .a(g849) );
  or2_316 OR2_271 ( .c(g11229), .b(g11154), .a(g11012) );
  or2_315 OR2_272 ( .c(g8973), .b(g8821), .a(g8735) );
  or2_314 OR2_273 ( .c(g10658), .b(g10595), .a(g7674) );
  or2_313 OR2_274 ( .c(g10339), .b(g10232), .a(g8574) );
  or4_40 OR4_21 ( .e(I5363), .d(g1149), .c(g1153), .b(g1157), .a(g1160) );
  or2_312 OR2_275 ( .c(g11310), .b(g11220), .a(g11100) );
  or2_311 OR2_276 ( .c(g6500), .b(g5725), .a(g4986) );
  or2_310 OR2_277 ( .c(g10855), .b(g6075), .a(g10736) );
  or2_309 OR2_278 ( .c(g9916), .b(g9855), .a(g9694) );
  or2_308 OR2_279 ( .c(g10411), .b(g10299), .a(g8574) );
  or2_307 OR2_280 ( .c(g11603), .b(g11582), .a(g11553) );
  or4_39 OR4_22 ( .e(I5357), .d(g1265), .c(g1260), .b(g1255), .a(g1250) );
  or2_306 OR2_281 ( .c(g9560), .b(g9052), .a(n1329) );
  or2_305 OR2_282 ( .c(g6672), .b(g4117), .a(g5259) );
  or3_39 OR3_23 ( .d(g9873), .c(g9623), .b(g9599), .a(g9758) );
  or2_304 OR2_283 ( .c(g6523), .b(g5745), .a(g4995) );
  or2_303 OR2_284 ( .c(g10707), .b(g5545), .a(g10686) );
  or4_38 OR4_23 ( .e(I5626), .d(g521), .c(g525), .b(g530), .a(g534) );
  or2_302 OR2_285 ( .c(g9579), .b(g9052), .a(n1329) );
  or2_301 OR2_286 ( .c(g7298), .b(g7136), .a(g6324) );
  or2_300 OR2_287 ( .c(g6551), .b(g5804), .a(g5031) );
  or2_299 OR2_288 ( .c(g6099), .b(g5273), .a(g4550) );
  or2_298 OR2_289 ( .c(g8282), .b(g8101), .a(g7819) );
  or2_297 OR2_290 ( .c(g9917), .b(g9856), .a(g9695) );
  or4_37 OR4_24 ( .e(I15057), .d(n1173), .c(g9680), .b(g9624), .a(g9785) );
  or2_296 OR2_291 ( .c(g7219), .b(g6661), .a(g4421) );
  or2_295 OR2_292 ( .c(g10019), .b(I15219), .a(I15220) );
  or2_294 OR2_293 ( .c(g5857), .b(g5418), .a(g4670) );
  or4_36 OR4_25 ( .e(g9725), .d(g9642), .c(g9659), .b(g9616), .a(I14862) );
  or2_293 OR2_294 ( .c(g11298), .b(g11212), .a(g11087) );
  or2_292 OR2_295 ( .c(g10402), .b(g10295), .a(g8574) );
  or4_35 OR4_26 ( .e(g2521), .d(g538), .c(g542), .b(g476), .a(I5626) );
  or3_38 OR3_24 ( .d(I14751), .c(g8995), .b(g9205), .a(g9192) );
  or2_291 OR2_296 ( .c(g10866), .b(g5539), .a(g10753) );
  or2_290 OR2_297 ( .c(g6534), .b(g5772), .a(g5003) );
  or2_289 OR2_298 ( .c(g11232), .b(g11158), .a(g11015) );
  or3_37 OR3_25 ( .d(g9706), .c(g9644), .b(g9386), .a(g9591) );
  or2_288 OR2_299 ( .c(g10001), .b(I15204), .a(I15205) );
  or2_287 OR2_300 ( .c(g8776), .b(g5510), .a(g8655) );
  or2_286 OR2_301 ( .c(g7225), .b(g6666), .a(g6079) );
  or3_36 OR3_26 ( .d(g9888), .c(g9648), .b(g9608), .a(g9757) );
  or2_285 OR2_302 ( .c(g11261), .b(g11238), .a(g11023) );
  or3_35 OR3_27 ( .d(g9956), .c(g9948), .b(g9942), .a(g9815) );
  or2_284 OR2_303 ( .c(g10923), .b(g10778), .a(g10715) );
  or2_283 OR2_304 ( .c(g8264), .b(g7879), .a(g3389) );
  or2_282 OR2_305 ( .c(g6513), .b(g5737), .a(g4991) );
  or3_34 OR3_28 ( .d(I14835), .c(g9621), .b(g9645), .a(g9588) );
  or2_281 OR2_306 ( .c(g8641), .b(g8120), .a(g8463) );
  or3_33 OR3_29 ( .d(g5361), .c(g4316), .b(n1392), .a(g126) );
  or2_280 OR2_307 ( .c(g11316), .b(g11226), .a(g11103) );
  or4_34 OR4_27 ( .e(I16161), .d(g10479), .c(g10478), .b(g10477), .a(g10475)
         );
  or2_279 OR2_308 ( .c(g6916), .b(g6348), .a(g5687) );
  or2_278 OR2_309 ( .c(g8777), .b(g5522), .a(g8659) );
  or4_33 OR4_28 ( .e(g2353), .d(g1403), .c(g1407), .b(g1411), .a(g1415) );
  or2_277 OR2_310 ( .c(g7510), .b(g7186), .a(g6730) );
  or3_32 OR3_30 ( .d(g9957), .c(g9949), .b(g9943), .a(g9776) );
  or2_276 OR2_311 ( .c(g2744), .b(I5804), .a(I5805) );
  or2_275 OR2_312 ( .c(g7245), .b(g6696), .a(g6102) );
  or2_274 OR2_313 ( .c(g7291), .b(g7050), .a(g6317) );
  or2_273 OR2_314 ( .c(g8611), .b(g8410), .a(g8556) );
  or4_32 OR4_29 ( .e(I15199), .d(g8167), .c(g9903), .b(g9932), .a(g9828) );
  or2_272 OR2_315 ( .c(g10550), .b(g1718), .a(g10450) );
  or2_271 OR2_316 ( .c(g11330), .b(g11304), .a(g11170) );
  or2_270 OR2_317 ( .c(g10721), .b(g10306), .a(g10669) );
  or2_269 OR2_318 ( .c(g8153), .b(g7888), .a(g6875) );
  or2_268 OR2_319 ( .c(g10773), .b(g5540), .a(g10685) );
  or2_267 OR2_320 ( .c(g3688), .b(n1392), .a(g868) );
  or4_31 OR4_30 ( .e(I15225), .d(g9842), .c(g9967), .b(g9859), .a(g9881) );
  or2_266 OR2_321 ( .c(g6042), .b(g5535), .a(g3987) );
  or2_265 OR2_322 ( .c(g10655), .b(g10561), .a(g7389) );
  or2_264 OR2_323 ( .c(g11259), .b(g11236), .a(g11021) );
  or2_263 OR2_324 ( .c(g11225), .b(g11149), .a(g11009) );
  or2_262 OR2_325 ( .c(g5914), .b(g5029), .a(g4343) );
  or2_261 OR2_326 ( .c(g11258), .b(g11235), .a(g11020) );
  or2_260 OR2_327 ( .c(g6054), .b(g5199), .a(g4483) );
  or3_31 OR3_31 ( .d(g9728), .c(g9412), .b(g9422), .a(g9426) );
  or3_30 OR3_32 ( .d(g9730), .c(g9414), .b(g9425), .a(g9423) );
  or2_259 OR2_328 ( .c(g5820), .b(g5595), .a(g4834) );
  or3_29 OR3_33 ( .d(g8574), .c(g30), .b(n1173), .a(n1184) );
  or2_258 OR2_329 ( .c(g11602), .b(g11581), .a(g11552) );
  or2_257 OR2_330 ( .c(g10502), .b(g4169), .a(g10365) );
  or2_256 OR2_331 ( .c(g10557), .b(g4123), .a(g10508) );
  or4_30 OR4_31 ( .e(I15171), .d(g8175), .c(g9909), .b(g9896), .a(g9835) );
  or2_255 OR2_332 ( .c(g11337), .b(g11282), .a(g11177) );
  or2_254 OR2_333 ( .c(g7465), .b(g6876), .a(g6410) );
  or2_253 OR2_334 ( .c(g8262), .b(g7970), .a(g7625) );
  or2_252 OR2_335 ( .c(g8889), .b(g8844), .a(g8756) );
  or2_251 OR2_336 ( .c(g7096), .b(g6544), .a(g5911) );
  or2_250 OR2_337 ( .c(g5995), .b(g5097), .a(g5099) );
  or2_249 OR2_338 ( .c(g8285), .b(g8104), .a(g7822) );
  or2_248 OR2_339 ( .c(g10791), .b(g6186), .a(g10762) );
  or2_247 OR2_340 ( .c(g2499), .b(I5570), .a(I5571) );
  or3_28 OR3_34 ( .d(I14607), .c(g8995), .b(g9205), .a(g9192) );
  or2_246 OR2_341 ( .c(g6049), .b(g5254), .a(g3718) );
  or2_245 OR2_342 ( .c(g9920), .b(g9860), .a(g9701) );
  or2_244 OR2_343 ( .c(g10556), .b(g4115), .a(g10506) );
  or2_243 OR2_344 ( .c(g8643), .b(g8364), .a(g8508) );
  or2_242 OR2_345 ( .c(g5810), .b(g5588), .a(g4823) );
  or2_241 OR2_346 ( .c(g11336), .b(g11281), .a(g11176) );
  or2_240 OR2_347 ( .c(g8742), .b(g8135), .a(g8598) );
  or2_239 OR2_348 ( .c(g8926), .b(g8848), .a(g8764) );
  or2_238 OR2_349 ( .c(g7218), .b(g6655), .a(g6070) );
  or4_29 OR4_32 ( .e(I15224), .d(g8174), .c(g9908), .b(g9937), .a(g9834) );
  or2_237 OR2_350 ( .c(g7293), .b(g7063), .a(g6319) );
  or2_236 OR2_351 ( .c(g11288), .b(g11204), .a(g11070) );
  or2_235 OR2_352 ( .c(g10800), .b(g6245), .a(g10772) );
  or2_234 OR2_353 ( .c(g11308), .b(g11218), .a(g11098) );
  or2_233 OR2_354 ( .c(g8269), .b(g7892), .a(g3429) );
  or2_232 OR2_355 ( .c(g10417), .b(g10301), .a(g8574) );
  or2_231 OR2_356 ( .c(g10936), .b(g5170), .a(g10808) );
  or2_230 OR2_357 ( .c(g9388), .b(n1330), .a(n1324) );
  or2_229 OR2_358 ( .c(g6185), .b(g5470), .a(g4715) );
  or2_228 OR2_359 ( .c(g6470), .b(g5699), .a(g4960) );
  or2_227 OR2_360 ( .c(g6897), .b(g6771), .a(g6240) );
  or2_226 OR2_361 ( .c(g8885), .b(g8841), .a(g8754) );
  or2_225 OR2_362 ( .c(g11260), .b(g11237), .a(g11022) );
  or2_224 OR2_363 ( .c(g11488), .b(g6671), .a(g11465) );
  or2_223 OR2_364 ( .c(g6105), .b(g5279), .a(g4559) );
  or2_222 OR2_365 ( .c(g10807), .b(g10701), .a(g10761) );
  or2_221 OR2_366 ( .c(g10639), .b(g10623), .a(g7734) );
  or2_220 OR2_367 ( .c(g4556), .b(g3536), .a(g1212) );
  or2_219 OR2_368 ( .c(g8288), .b(g8119), .a(g7825) );
  or2_218 OR2_369 ( .c(g6755), .b(g3524), .a(g5479) );
  or3_27 OR3_35 ( .d(I14862), .c(g9587), .b(g9600), .a(g9611) );
  or4_28 OR4_33 ( .e(I16160), .d(g10394), .c(g10392), .b(g10482), .a(g10481)
         );
  or4_27 OR4_34 ( .e(I15042), .d(n1173), .c(g9686), .b(g9624), .a(g9785) );
  or2_217 OR2_370 ( .c(g11610), .b(g11589), .a(g11560) );
  or4_26 OR4_35 ( .e(g9711), .d(g9660), .c(g9390), .b(g9359), .a(g9589) );
  or2_216 OR2_371 ( .c(g6045), .b(g5541), .a(g3989) );
  or2_215 OR2_372 ( .c(g11270), .b(g11198), .a(g11032) );
  or2_214 OR2_373 ( .c(g7258), .b(g6549), .a(g5913) );
  or2_213 OR2_374 ( .c(g6059), .b(g5211), .a(g4489) );
  or2_212 OR2_375 ( .c(g10007), .b(I15209), .a(I15210) );
  or2_211 OR2_376 ( .c(g11267), .b(g11192), .a(g11029) );
  or2_210 OR2_377 ( .c(g11294), .b(g6576), .a(g11210) );
  or3_26 OR3_36 ( .d(g9509), .c(n1325), .b(g9125), .a(g9111) );
  or2_209 OR2_378 ( .c(g7211), .b(g6647), .a(g6067) );
  or2_208 OR2_379 ( .c(g5404), .b(g4487), .a(g3696) );
  or2_207 OR2_380 ( .c(g4089), .b(g1959), .a(n1302) );
  or4_25 OR4_36 ( .e(I15219), .d(g8172), .c(g9907), .b(g9936), .a(g9833) );
  or2_206 OR2_381 ( .c(g11219), .b(g11145), .a(g11006) );
  or2_205 OR2_382 ( .c(g6015), .b(g5497), .a(g3942) );
  or2_204 OR2_383 ( .c(g10720), .b(g10304), .a(g10667) );
  or2_203 OR2_384 ( .c(g8265), .b(g7881), .a(g3396) );
  or2_202 OR2_385 ( .c(g5224), .b(g4360), .a(g3512) );
  or3_25 OR3_37 ( .d(g9700), .c(g9358), .b(g9667), .a(I14827) );
  or2_201 OR2_386 ( .c(g7106), .b(g6554), .a(g5917) );
  or2_200 OR2_387 ( .c(g8770), .b(g5476), .a(g8651) );
  or2_199 OR2_388 ( .c(g11201), .b(g11152), .a(g11011) );
  or3_24 OR3_38 ( .d(g9950), .c(g9901), .b(g9898), .a(g9779) );
  or4_24 OR4_37 ( .e(g9723), .d(g9620), .c(g9652), .b(g9391), .a(I14858) );
  or2_198 OR2_389 ( .c(g2309), .b(I5357), .a(I5358) );
  or2_197 OR2_390 ( .c(g11266), .b(g11190), .a(g11028) );
  or2_196 OR2_391 ( .c(g10727), .b(g4969), .a(g10638) );
  or2_195 OR2_392 ( .c(g10863), .b(g5531), .a(g10750) );
  or2_194 OR2_393 ( .c(g8429), .b(g8385), .a(g8069) );
  or2_193 OR2_394 ( .c(g9751), .b(g9515), .a(g9510) );
  or2_192 OR2_395 ( .c(g8281), .b(g8097), .a(g7818) );
  or2_191 OR2_396 ( .c(g6910), .b(g6341), .a(g5680) );
  or2_190 OR2_397 ( .c(g8639), .b(g8118), .a(g8462) );
  or3_23 OR3_39 ( .d(g9673), .c(n1327), .b(n1331), .a(n1323) );
  or2_189 OR2_398 ( .c(g11285), .b(g11255), .a(g11161) );
  or2_188 OR2_399 ( .c(g11305), .b(g11215), .a(g11093) );
  or4_23 OR4_38 ( .e(I15177), .d(g9844), .c(g9960), .b(g9863), .a(g9876) );
  or3_22 OR3_40 ( .d(g9734), .c(g9415), .b(g9428), .a(g9421) );
  or3_21 OR3_41 ( .d(I14827), .c(g9603), .b(g9614), .a(g9584) );
  or2_187 OR2_400 ( .c(g5824), .b(g5602), .a(g4839) );
  or2_186 OR2_401 ( .c(g8715), .b(g8416), .a(g8687) );
  or2_185 OR2_402 ( .c(g5762), .b(g5178), .a(g5186) );
  or2_184 OR2_403 ( .c(g6538), .b(g5782), .a(g5006) );
  or2_183 OR2_404 ( .c(g5590), .b(g4718), .a(g4723) );
  or2_182 OR2_405 ( .c(g10726), .b(g10316), .a(g10673) );
  or2_181 OR2_406 ( .c(g3120), .b(I6350), .a(I6351) );
  or2_180 OR2_407 ( .c(g9573), .b(g9052), .a(n1329) );
  or3_20 OR3_42 ( .d(g4640), .c(n1392), .b(g3563), .a(g1527) );
  or2_179 OR2_408 ( .c(g6093), .b(g5264), .a(g4534) );
  or2_178 OR2_409 ( .c(g8162), .b(g7898), .a(g6889) );
  or2_177 OR2_410 ( .c(g8268), .b(g7962), .a(g7613) );
  or2_176 OR2_411 ( .c(g9569), .b(g9052), .a(n1329) );
  or2_175 OR2_412 ( .c(g11485), .b(g6646), .a(g11462) );
  or2_174 OR2_413 ( .c(g10797), .b(g6206), .a(g10766) );
  or3_19 OR3_43 ( .d(I14779), .c(g8995), .b(g9205), .a(g9192) );
  or2_173 OR2_414 ( .c(g10408), .b(g10298), .a(g8574) );
  or2_172 OR2_415 ( .c(g10635), .b(g10622), .a(g7732) );
  or2_171 OR2_416 ( .c(g2305), .b(I5351), .a(I5352) );
  or4_22 OR4_39 ( .e(I15176), .d(g8176), .c(g9910), .b(g9897), .a(g9836) );
  or2_170 OR2_417 ( .c(g3435), .b(g2945), .a(g2950) );
  or2_169 OR2_418 ( .c(g9924), .b(g9866), .a(g9709) );
  or2_168 OR2_419 ( .c(g10711), .b(g5547), .a(g10690) );
  or2_167 OR2_420 ( .c(g5814), .b(g5591), .a(g4827) );
  or2_166 OR2_421 ( .c(g5038), .b(g4878), .a(g4884) );
  or4_21 OR4_40 ( .e(I15215), .d(g9840), .c(g9965), .b(g9854), .a(g9879) );
  or2_165 OR2_422 ( .c(g8226), .b(g7504), .a(g82) );
  or2_164 OR2_423 ( .c(g7367), .b(g7224), .a(g6744) );
  or2_163 OR2_424 ( .c(g7457), .b(g6873), .a(g6404) );
  or2_162 OR2_425 ( .c(g5229), .b(g4364), .a(g3516) );
  or2_161 OR2_426 ( .c(g5993), .b(g5090), .a(g4400) );
  or2_160 OR2_427 ( .c(g8283), .b(g8098), .a(g7820) );
  or2_159 OR2_428 ( .c(g7971), .b(g5110), .a(g7549) );
  or2_158 OR2_429 ( .c(g8602), .b(g8401), .a(g8550) );
  or2_157 OR2_430 ( .c(g8920), .b(g8845), .a(g8759) );
  or2_156 OR2_431 ( .c(g10663), .b(g10237), .a(g10581) );
  or2_155 OR2_432 ( .c(g6074), .b(g5349), .a(g1) );
  or2_154 OR2_433 ( .c(g8261), .b(g7876), .a(g3383) );
  or2_153 OR2_434 ( .c(g10862), .b(g5524), .a(g10746) );
  or2_152 OR2_435 ( .c(g5837), .b(g5640), .a(g4224) );
  or2_151 OR2_436 ( .c(g11333), .b(g11274), .a(g11173) );
  or2_150 OR2_437 ( .c(g6080), .b(g5249), .a(g4512) );
  or2_149 OR2_438 ( .c(g6480), .b(g5721), .a(g4971) );
  or2_148 OR2_439 ( .c(g7740), .b(g7209), .a(g6741) );
  or2_147 OR2_440 ( .c(g10702), .b(g10562), .a(g2984) );
  or3_18 OR3_44 ( .d(g9697), .c(g9665), .b(g9606), .a(I14822) );
  or2_146 OR2_441 ( .c(g8203), .b(g7453), .a(n1383) );
  or2_145 OR2_442 ( .c(g9914), .b(g9851), .a(g9692) );
  or2_144 OR2_443 ( .c(g10564), .b(g10560), .a(g7368) );
  or2_143 OR2_444 ( .c(g11484), .b(g6639), .a(g11461) );
  or2_142 OR2_445 ( .c(g5842), .b(g5618), .a(g4870) );
  or4_20 OR4_41 ( .e(I15200), .d(g9837), .c(g9962), .b(g9848), .a(g9880) );
  or2_141 OR2_446 ( .c(g11609), .b(g11588), .a(g11559) );
  or3_17 OR3_45 ( .d(I14582), .c(g8995), .b(g9205), .a(g9192) );
  or2_140 OR2_447 ( .c(g8940), .b(g8793), .a(g8703) );
  or2_139 OR2_448 ( .c(g11312), .b(g11222), .a(g11101) );
  or2_138 OR2_449 ( .c(g11608), .b(g11587), .a(g11558) );
  or2_137 OR2_450 ( .c(g6000), .b(g5480), .a(g3912) );
  or2_136 OR2_451 ( .c(g8428), .b(g8382), .a(g8068) );
  or2_135 OR2_452 ( .c(g8430), .b(g8386), .a(g8070) );
  or2_134 OR2_453 ( .c(g9922), .b(g9864), .a(g9705) );
  or2_133 OR2_454 ( .c(g8247), .b(g8010), .a(g7704) );
  or2_132 OR2_455 ( .c(g3438), .b(g2939), .a(g2944) );
  or4_19 OR4_42 ( .e(I5576), .d(g431), .c(g435), .b(g440), .a(g444) );
  or2_131 OR2_456 ( .c(g6924), .b(g6362), .a(g4261) );
  or2_130 OR2_457 ( .c(g5405), .b(g4476), .a(n1264) );
  or2_129 OR2_458 ( .c(g8638), .b(g8108), .a(g8461) );
  or2_128 OR2_459 ( .c(g8609), .b(g8408), .a(g8555) );
  or2_127 OR2_460 ( .c(g9995), .b(I15199), .a(I15200) );
  or2_126 OR2_461 ( .c(g8883), .b(g8838), .a(g8753) );
  or4_18 OR4_43 ( .e(I15214), .d(g8170), .c(g9906), .b(g9935), .a(g9831) );
  or3_16 OR3_46 ( .d(g2538), .c(g1466), .b(g1458), .a(I5649) );
  or2_125 OR2_462 ( .c(g11329), .b(g11302), .a(g11169) );
  or2_124 OR2_463 ( .c(g4255), .b(g4009), .a(g4047) );
  or2_123 OR2_464 ( .c(g11328), .b(g11299), .a(g11168) );
  or3_15 OR3_47 ( .d(g9704), .c(g9385), .b(g9605), .a(I14835) );
  or4_17 OR4_44 ( .e(I5352), .d(g1129), .c(g1125), .b(g1121), .a(g1117) );
  or2_122 OR2_465 ( .c(g8774), .b(g5499), .a(g8654) );
  or3_14 OR3_48 ( .d(g9954), .c(g9946), .b(g9940), .a(g9781) );
  or2_121 OR2_466 ( .c(g10405), .b(g10297), .a(g8574) );
  or2_120 OR2_467 ( .c(g9363), .b(g9205), .a(g9192) );
  or2_119 OR2_468 ( .c(g5849), .b(g4949), .a(g4144) );
  or4_16 OR4_45 ( .e(I5599), .d(g516), .c(g511), .b(g506), .a(g501) );
  or2_118 OR2_469 ( .c(g7204), .b(g6645), .a(g4421) );
  or2_117 OR2_470 ( .c(g7300), .b(g7139), .a(g6326) );
  or2_116 OR2_471 ( .c(g4293), .b(g4064), .a(g4068) );
  or2_115 OR2_472 ( .c(g9912), .b(g9847), .a(g9690) );
  or2_114 OR2_473 ( .c(g6533), .b(g5771), .a(g5002) );
  or2_113 OR2_474 ( .c(g8816), .b(g7951), .a(g8731) );
  or2_112 OR2_475 ( .c(g9929), .b(g9871), .a(g9718) );
  or2_111 OR2_476 ( .c(g5819), .b(g5625), .a(g4876) );
  or3_13 OR3_49 ( .d(I14831), .c(g9613), .b(g9622), .a(g9586) );
  or2_110 OR2_477 ( .c(g5852), .b(g5632), .a(g4883) );
  or2_109 OR2_478 ( .c(g8263), .b(g8032), .a(g7720) );
  or2_108 OR2_479 ( .c(g3431), .b(g2951), .a(g2957) );
  or3_12 OR3_50 ( .d(g9683), .c(n1327), .b(n1331), .a(n1323) );
  or2_107 OR2_480 ( .c(g8631), .b(g8474), .a(g7449) );
  or2_106 OR2_481 ( .c(g6922), .b(g6352), .a(g5694) );
  or2_105 OR2_482 ( .c(g8817), .b(g7954), .a(g8732) );
  or4_15 OR4_46 ( .e(g9735), .d(g9649), .c(g9651), .b(g9384), .a(g9361) );
  or2_104 OR2_483 ( .c(g8605), .b(g8404), .a(g8553) );
  or2_103 OR2_484 ( .c(g11263), .b(g11187), .a(g11025) );
  or2_102 OR2_485 ( .c(g6739), .b(g5769), .a(g5780) );
  or2_101 OR2_486 ( .c(g11332), .b(g11273), .a(g11172) );
  or2_100 OR2_487 ( .c(g7143), .b(g6619), .a(g4421) );
  or2_99 OR2_488 ( .c(g6479), .b(g5707), .a(g4968) );
  or4_14 OR4_47 ( .e(I15048), .d(n1173), .c(g9683), .b(g9624), .a(g9785) );
  or2_98 OR2_489 ( .c(g6501), .b(g5726), .a(g4987) );
  or3_11 OR3_51 ( .d(g9702), .c(g9365), .b(g9647), .a(I14831) );
  or2_97 OR2_490 ( .c(g11221), .b(g11146), .a(g11007) );
  or3_10 OR3_52 ( .d(g9952), .c(g9944), .b(g9938), .a(g9817) );
  or2_96 OR2_491 ( .c(g11613), .b(g11600), .a(g11591) );
  or2_95 OR2_492 ( .c(g7621), .b(g5108), .a(g6994) );
  or2_94 OR2_493 ( .c(g3399), .b(g2918), .a(g2940) );
  or2_93 OR2_494 ( .c(g11605), .b(g11584), .a(g11555) );
  or2_92 OR2_495 ( .c(g4274), .b(g4054), .a(g4058) );
  or3_9 OR3_53 ( .d(I14602), .c(g8995), .b(g9205), .a(g9192) );
  or4_13 OR4_48 ( .e(I15033), .d(n1173), .c(n1327), .b(g9624), .a(g9785) );
  or2_91 OR2_496 ( .c(g10717), .b(g6235), .a(g10705) );
  or3_8 OR3_54 ( .d(I5629), .c(g845), .b(g841), .a(g837) );
  or2_90 OR2_497 ( .c(g9925), .b(g9867), .a(g9712) );
  or2_89 OR2_498 ( .c(g3819), .b(g3275), .a(g9) );
  or2_88 OR2_499 ( .c(g6912), .b(g6350), .a(g4235) );
  or2_87 OR2_500 ( .c(g10723), .b(g4952), .a(g10633) );
  or2_86 OR2_501 ( .c(g6929), .b(g6360), .a(g5704) );
  or2_85 OR2_502 ( .c(g10646), .b(g10625), .a(g7739) );
  or2_84 OR2_503 ( .c(g9516), .b(n1325), .a(g9125) );
  or2_83 OR2_504 ( .c(g6626), .b(g5934), .a(g123) );
  or4_12 OR4_49 ( .e(I6350), .d(g2445), .c(g2437), .b(g2433), .a(g2419) );
  or2_82 OR2_505 ( .c(g11325), .b(g11295), .a(g11165) );
  or4_11 OR4_50 ( .e(I5366), .d(g1280), .c(g1284), .b(g1292), .a(g1296) );
  or3_7 OR3_55 ( .d(I5649), .c(g1499), .b(g1486), .a(g1482) );
  or2_81 OR2_506 ( .c(g6894), .b(g6763), .a(g4868) );
  or3_6 OR3_56 ( .d(g9738), .c(g9417), .b(g9447), .a(g9506) );
  or2_80 OR2_507 ( .c(g8383), .b(g8163), .a(g5051) );
  or2_79 OR2_508 ( .c(g8779), .b(g5530), .a(g8663) );
  or2_78 OR2_509 ( .c(g8161), .b(g8005), .a(g7185) );
  or2_77 OR2_510 ( .c(g8451), .b(n1264), .a(g8366) );
  or2_76 OR2_511 ( .c(g9915), .b(g9853), .a(g9693) );
  or4_10 OR4_51 ( .e(g2316), .d(g1300), .c(g1304), .b(g1270), .a(I5366) );
  or2_75 OR2_512 ( .c(g5576), .b(g4675), .a(n1254) );
  or2_74 OR2_513 ( .c(g10857), .b(g6090), .a(g10738) );
  or2_73 OR2_514 ( .c(g10793), .b(g6194), .a(g10763) );
  or2_72 OR2_515 ( .c(g7511), .b(g6890), .a(g6438) );
  or2_71 OR2_516 ( .c(g8944), .b(g8799), .a(g8708) );
  or2_70 OR2_517 ( .c(g10765), .b(g5492), .a(g10680) );
  or2_69 OR2_518 ( .c(g10549), .b(g1718), .a(g10451) );
  or2_68 OR2_519 ( .c(g7092), .b(g6540), .a(g5902) );
  or2_67 OR2_520 ( .c(g11604), .b(g11583), .a(g11554) );
  or2_66 OR2_521 ( .c(g8434), .b(g8400), .a(g8074) );
  or2_65 OR2_522 ( .c(g6546), .b(g5796), .a(g5026) );
  or2_64 OR2_523 ( .c(g3354), .b(n1392), .a(g1216) );
  or2_63 OR2_524 ( .c(g9928), .b(g9870), .a(g9717) );
  or2_62 OR2_525 ( .c(g11262), .b(g11240), .a(g11024) );
  or4_9 OR4_52 ( .e(g9785), .d(n1326), .c(g8995), .b(g9388), .a(g9363) );
  or2_61 OR2_526 ( .c(g5867), .b(n1264), .a(g4921) );
  or2_60 OR2_527 ( .c(g8210), .b(g7466), .a(n1383) );
  or2_59 OR2_528 ( .c(g10533), .b(g1718), .a(g10449) );
  or2_58 OR2_529 ( .c(g9563), .b(g9052), .a(n1329) );
  or2_57 OR2_530 ( .c(g6906), .b(g6791), .a(g5674) );
  or2_56 OR2_531 ( .c(g7375), .b(g7230), .a(g6745) );
  or2_55 OR2_532 ( .c(g7651), .b(g7135), .a(n1392) );
  or4_8 OR4_53 ( .e(I5570), .d(g416), .c(g411), .b(g406), .a(g401) );
  or3_5 OR3_57 ( .d(g9731), .c(g9641), .b(g9364), .a(g9387) );
  or2_54 OR2_533 ( .c(g11247), .b(g11097), .a(g10949) );
  or4_7 OR4_54 ( .e(I15045), .d(n1173), .c(g9676), .b(g9624), .a(g9785) );
  or2_53 OR2_534 ( .c(g10856), .b(g6083), .a(g10737) );
  or2_52 OR2_535 ( .c(g9557), .b(g9052), .a(n1329) );
  or2_51 OR2_536 ( .c(g7184), .b(g6625), .a(g6047) );
  or2_50 OR2_537 ( .c(g11612), .b(g11599), .a(g11590) );
  or2_49 OR2_538 ( .c(g7384), .b(g7088), .a(g6618) );
  or2_48 OR2_539 ( .c(g11324), .b(g11271), .a(g11164) );
  or2_47 OR2_540 ( .c(g8922), .b(g8822), .a(g8736) );
  or4_6 OR4_55 ( .e(I5358), .d(g1245), .c(g1240), .b(g1235), .a(g1275) );
  or3_4 OR3_58 ( .d(g9955), .c(g9947), .b(g9941), .a(g9808) );
  or4_5 OR4_56 ( .e(g2501), .d(g448), .c(g452), .b(g421), .a(I5576) );
  or2_46 OR2_541 ( .c(g7231), .b(g6673), .a(g6087) );
  or2_45 OR2_542 ( .c(g6078), .b(g4503), .a(g5256) );
  or2_44 OR2_543 ( .c(g6478), .b(g5706), .a(g4967) );
  or2_43 OR2_544 ( .c(g6907), .b(g6792), .a(g5675) );
  or2_42 OR2_545 ( .c(g6035), .b(g5518), .a(g3974) );
  or2_41 OR2_546 ( .c(g8937), .b(g8786), .a(g8698) );
  or2_40 OR2_547 ( .c(g7742), .b(g7217), .a(g6743) );
  or2_39 OR2_548 ( .c(g10722), .b(g10308), .a(g10671) );
  or2_38 OR2_549 ( .c(g9918), .b(g9858), .a(g9698) );
  or2_37 OR2_550 ( .c(g5403), .b(g4486), .a(g3695) );
  or2_36 OR2_551 ( .c(g7926), .b(g7435), .a(g6892) );
  or2_35 OR2_552 ( .c(g6915), .b(g6347), .a(g5686) );
  or2_34 OR2_553 ( .c(g5841), .b(g4914), .a(g4230) );
  or4_4 OR4_57 ( .e(I15220), .d(g9841), .c(g9966), .b(g9857), .a(g9877) );
  or2_33 OR2_554 ( .c(g10529), .b(I16160), .a(I16161) );
  or2_32 OR2_555 ( .c(g11246), .b(g11094), .a(g10948) );
  or2_31 OR2_556 ( .c(g6002), .b(g5489), .a(g3939) );
  or2_30 OR2_557 ( .c(g7712), .b(g7125), .a(n1392) );
  or2_29 OR2_558 ( .c(g8810), .b(g7933), .a(g8720) );
  or2_28 OR2_559 ( .c(g9921), .b(g9862), .a(g9703) );
  or2_27 OR2_560 ( .c(g8432), .b(g8389), .a(g8072) );
  or4_3 OR4_58 ( .e(I15172), .d(g9843), .c(g9959), .b(g9861), .a(g9874) );
  or3_3 OR3_59 ( .d(I14822), .c(g9597), .b(g9604), .a(g9582) );
  or2_26 OR2_561 ( .c(g6928), .b(g6359), .a(g5703) );
  or2_25 OR2_562 ( .c(g8157), .b(n1245), .a(g7623) );
  or2_24 OR2_563 ( .c(g6930), .b(g6364), .a(g4269) );
  or2_23 OR2_564 ( .c(g7660), .b(g7059), .a(g5867) );
  or2_22 OR2_565 ( .c(g6899), .b(g6463), .a(g32) );
  or2_21 OR2_566 ( .c(g9392), .b(g9328), .a(g9324) );
  or2_20 OR2_567 ( .c(g11318), .b(g11228), .a(g11104) );
  or3_2 OR3_60 ( .d(I16427), .c(n1297), .b(g10383), .a(g10382) );
  or2_19 OR2_568 ( .c(g11227), .b(g11151), .a(g11010) );
  or2_18 OR2_569 ( .c(g11058), .b(g10933), .a(g5280) );
  or4_2 OR4_59 ( .e(I5351), .d(g1145), .c(g1141), .b(g1137), .a(g1133) );
  or3_1 OR3_61 ( .d(g9708), .c(g9653), .b(g9389), .a(g9646) );
  or2_17 OR2_570 ( .c(g6071), .b(g5228), .a(g4505) );
  or2_16 OR2_571 ( .c(g9911), .b(g9846), .a(g9689) );
  or2_15 OR2_572 ( .c(g7102), .b(g6550), .a(g5915) );
  or2_14 OR2_573 ( .c(g7302), .b(g7141), .a(g6328) );
  or2_13 OR2_574 ( .c(g6038), .b(g5528), .a(g3979) );
  or2_12 OR2_575 ( .c(g4239), .b(g4000), .a(g4008) );
  or2_11 OR2_576 ( .c(g8646), .b(g8224), .a(g8547) );
  or2_10 OR2_577 ( .c(g9974), .b(I15176), .a(I15177) );
  or2_9 OR2_578 ( .c(g5823), .b(g5631), .a(g4882) );
  or2_8 OR2_579 ( .c(g6918), .b(g6358), .a(g4252) );
  or2_7 OR2_580 ( .c(g7265), .b(g6756), .a(g6204) );
  or4_1 OR4_60 ( .e(I5804), .d(g2111), .c(g2109), .b(g2106), .a(g2104) );
  or2_6 OR2_581 ( .c(g5851), .b(g4941), .a(g4253) );
  or2_5 OR2_582 ( .c(g11481), .b(g6624), .a(g11458) );
  or2_4 OR2_583 ( .c(g10336), .b(g10230), .a(g8574) );
  or2_3 OR2_584 ( .c(g7296), .b(g7131), .a(g6322) );
  or2_2 OR2_585 ( .c(g4300), .b(n1392), .a(g1212) );
  or2_1 OR2_586 ( .c(g8647), .b(g8130), .a(g8470) );
  nand2_0 NAND2_0 ( .c(g8546), .b(n1278), .a(g8390) );
  nand2_923 NAND2_1 ( .c(g2516), .b(I5612), .a(I5613) );
  nand2_922 NAND2_2 ( .c(g2987), .b(n1072), .a(g883) );
  nand2_921 NAND2_3 ( .c(I5593), .b(g1703), .a(I5591) );
  nand2_920 NAND2_4 ( .c(g8970), .b(g5548), .a(g8839) );
  nand2_919 NAND2_5 ( .c(I10519), .b(g6231), .a(g822) );
  nand2_918 NAND2_6 ( .c(I11279), .b(g305), .a(I11278) );
  nand4_0 NAND4_0 ( .e(g7990), .d(n1311), .c(n1310), .b(g43), .a(g42) );
  nand2_917 NAND2_7 ( .c(I11278), .b(g305), .a(g6485) );
  nand2_916 NAND2_8 ( .c(g3978), .b(n1289), .a(g1822) );
  nand2_915 NAND2_9 ( .c(I5264), .b(n1336), .a(I5263) );
  nand2_914 NAND2_10 ( .c(I8640), .b(g4278), .a(g516) );
  nand2_913 NAND2_11 ( .c(I6761), .b(g2943), .a(I6760) );
  nand2_912 NAND2_12 ( .c(I17400), .b(g11418), .a(g11416) );
  nand2_911 NAND2_13 ( .c(I5450), .b(g1235), .a(I5449) );
  nand2_910 NAND2_14 ( .c(I16060), .b(g10372), .a(I16058) );
  nand2_909 NAND2_15 ( .c(I6746), .b(g2938), .a(g1453) );
  nand2_908 NAND2_16 ( .c(I11975), .b(g1462), .a(I11973) );
  nand2_907 NAND2_17 ( .c(I12136), .b(g6038), .a(g131) );
  nand2_906 NAND2_18 ( .c(I11937), .b(g1458), .a(I11935) );
  nand2_905 NAND2_19 ( .c(g2959), .b(I6167), .a(I6168) );
  nand2_904 NAND2_20 ( .c(I5878), .b(g2120), .a(g2115) );
  nand2_903 NAND2_21 ( .c(g2517), .b(I5619), .a(I5620) );
  nand2_902 NAND2_22 ( .c(g5552), .b(n1265), .a(g4401) );
  nand2_901 NAND2_23 ( .c(I6468), .b(g23), .a(I6467) );
  nand2_900 NAND2_24 ( .c(I8796), .b(g4672), .a(I8795) );
  nand2_899 NAND2_25 ( .c(g10392), .b(I15891), .a(I15892) );
  nand2_898 NAND2_26 ( .c(I5611), .b(g1280), .a(g1284) );
  nand2_897 NAND2_27 ( .c(g8738), .b(n1261), .a(g4921) );
  nand2_896 NAND2_28 ( .c(I6716), .b(g201), .a(I6714) );
  nand2_895 NAND2_29 ( .c(g2310), .b(g591), .a(g605) );
  nand2_894 NAND2_30 ( .c(I7685), .b(g3460), .a(I7683) );
  nand2_893 NAND2_31 ( .c(g3056), .b(n1126), .a(g599) );
  nand2_892 NAND2_32 ( .c(I12108), .b(g135), .a(I12106) );
  nand3_0 NAND3_0 ( .d(g3529), .c(g2310), .b(g3062), .a(g2325) );
  nand2_891 NAND2_33 ( .c(I6747), .b(g2938), .a(I6746) );
  nand2_890 NAND2_34 ( .c(g2236), .b(I5230), .a(I5231) );
  nand2_889 NAND2_35 ( .c(g7584), .b(I12075), .a(I12076) );
  nand2_888 NAND2_36 ( .c(I15870), .b(g10358), .a(g1796) );
  nand2_887 NAND2_37 ( .c(I16067), .b(g1806), .a(I16065) );
  nand2_886 NAND2_38 ( .c(I7562), .b(g3533), .a(g654) );
  nand2_885 NAND2_39 ( .c(I13531), .b(g8253), .a(I13529) );
  nand2_884 NAND2_40 ( .c(I8797), .b(g1145), .a(I8795) );
  nand2_883 NAND2_41 ( .c(I17584), .b(g11217), .a(n1293) );
  nand2_882 NAND2_42 ( .c(I11936), .b(g5857), .a(I11935) );
  nand2_881 NAND2_43 ( .c(I15257), .b(g9974), .a(I15256) );
  nand2_880 NAND2_44 ( .c(g8402), .b(I13505), .a(I13506) );
  nand3_22 NAND3_1 ( .d(g8824), .c(g8502), .b(g8501), .a(g8512) );
  nand2_879 NAND2_45 ( .c(I6186), .b(g2511), .a(n1335) );
  nand2_878 NAND2_46 ( .c(g11496), .b(I17504), .a(I17505) );
  nand2_877 NAND2_47 ( .c(I16001), .b(g1771), .a(I15999) );
  nand2_876 NAND2_48 ( .c(I6125), .b(g2215), .a(I6124) );
  nand2_875 NAND2_49 ( .c(I11909), .b(g1474), .a(I11907) );
  nand2_874 NAND2_50 ( .c(I12040), .b(g1466), .a(I12038) );
  nand2_873 NAND2_51 ( .c(I13909), .b(g1432), .a(I13907) );
  nand2_872 NAND2_52 ( .c(g3625), .b(I6771), .a(I6772) );
  nand2_871 NAND2_53 ( .c(I11908), .b(g5838), .a(I11907) );
  nand2_870 NAND2_54 ( .c(g10470), .b(I16008), .a(I16009) );
  nand2_869 NAND2_55 ( .c(I13908), .b(g8265), .a(I13907) );
  nand2_868 NAND2_56 ( .c(g3813), .b(I7034), .a(I7035) );
  nand2_867 NAND2_57 ( .c(I8650), .b(g4824), .a(g778) );
  nand2_866 NAND2_58 ( .c(g6207), .b(I9947), .a(I9948) );
  nand2_865 NAND2_59 ( .c(I16066), .b(g10428), .a(I16065) );
  nand2_864 NAND2_60 ( .c(g2948), .b(I6144), .a(I6145) );
  nand2_863 NAND2_61 ( .c(I11242), .b(g6760), .a(I11241) );
  nand2_862 NAND2_62 ( .c(g10467), .b(I15993), .a(I15994) );
  nand2_861 NAND2_63 ( .c(I6187), .b(g2511), .a(I6186) );
  nand2_860 NAND2_64 ( .c(g6488), .b(g6027), .a(g6019) );
  nand2_859 NAND2_65 ( .c(I5500), .b(g1255), .a(g1007) );
  nand2_858 NAND2_66 ( .c(I11974), .b(g5852), .a(I11973) );
  nand2_857 NAND2_67 ( .c(I12062), .b(g1478), .a(I12060) );
  nand2_856 NAND2_68 ( .c(g5300), .b(I8771), .a(I8772) );
  nand2_855 NAND2_69 ( .c(I5184), .b(g1415), .a(g1515) );
  nand2_854 NAND2_70 ( .c(I13293), .b(g1882), .a(g8161) );
  nand2_853 NAND2_71 ( .c(I6200), .b(g2525), .a(I6199) );
  nand2_852 NAND2_72 ( .c(I13265), .b(g1909), .a(g8154) );
  nand2_851 NAND2_73 ( .c(I5024), .b(g995), .a(I5023) );
  nand2_850 NAND2_74 ( .c(I7863), .b(g4099), .a(g774) );
  nand2_849 NAND2_75 ( .c(g8705), .b(I13991), .a(I13992) );
  nand2_848 NAND2_76 ( .c(g8471), .b(I13660), .a(I13661) );
  nand2_847 NAND2_77 ( .c(I15256), .b(g9974), .a(g9968) );
  nand2_846 NAND2_78 ( .c(I6145), .b(g646), .a(I6143) );
  nand2_845 NAND2_79 ( .c(I13992), .b(n1261), .a(I13990) );
  nand2_844 NAND2_80 ( .c(I11510), .b(g1806), .a(I11508) );
  nand2_843 NAND2_81 ( .c(g10853), .b(g10731), .a(g5034) );
  nand2_842 NAND2_82 ( .c(I5231), .b(g148), .a(I5229) );
  nand2_841 NAND2_83 ( .c(I12047), .b(g1486), .a(I12045) );
  nand2_840 NAND2_84 ( .c(I10771), .b(g1801), .a(I10769) );
  nand2_839 NAND2_85 ( .c(g10477), .b(I16045), .a(I16046) );
  nand2_838 NAND2_86 ( .c(g7582), .b(I12061), .a(I12062) );
  nand2_837 NAND2_87 ( .c(I5104), .b(g431), .a(g435) );
  nand2_836 NAND2_88 ( .c(g8409), .b(I13530), .a(I13531) );
  nand2_835 NAND2_89 ( .c(I6447), .b(g2264), .a(g1776) );
  nand2_834 NAND2_90 ( .c(I4956), .b(g327), .a(I4954) );
  nand2_833 NAND2_91 ( .c(I5613), .b(g1284), .a(I5611) );
  nand2_832 NAND2_92 ( .c(I8481), .b(g3530), .a(I8479) );
  nand2_831 NAND2_93 ( .c(g5278), .b(I8739), .a(I8740) );
  nand2_830 NAND2_94 ( .c(I6880), .b(g3301), .a(I6879) );
  nand2_829 NAND2_95 ( .c(I15431), .b(g10001), .a(I15430) );
  nand2_828 NAND2_96 ( .c(g5548), .b(g1840), .a(g4401) );
  nand4_20 NAND4_1 ( .e(g7671), .d(n1311), .c(n1310), .b(n1309), .a(n1308) );
  nand2_827 NAND2_97 ( .c(I12020), .b(g6049), .a(I12019) );
  nand2_826 NAND2_98 ( .c(g10665), .b(I16331), .a(I16332) );
  nand2_825 NAND2_99 ( .c(I16469), .b(g10518), .a(I16467) );
  nand2_824 NAND2_100 ( .c(I5014), .b(g1007), .a(I5013) );
  nand2_823 NAND2_101 ( .c(I13523), .b(g8249), .a(I13521) );
  nand2_822 NAND2_102 ( .c(I16039), .b(g1791), .a(I16037) );
  nand2_821 NAND2_103 ( .c(I16468), .b(g10716), .a(I16467) );
  nand2_820 NAND2_104 ( .c(I12046), .b(g5814), .a(I12045) );
  nand2_819 NAND2_105 ( .c(g4476), .b(g3807), .a(g3071) );
  nand2_818 NAND2_106 ( .c(g10476), .b(I16038), .a(I16039) );
  nand2_817 NAND2_107 ( .c(I16038), .b(g10427), .a(I16037) );
  nand2_816 NAND2_108 ( .c(I8676), .b(g4374), .a(g1027) );
  nand2_815 NAND2_109 ( .c(I12113), .b(g6002), .a(g162) );
  nand2_814 NAND2_110 ( .c(I8761), .b(g4616), .a(g1129) );
  nand2_813 NAND2_111 ( .c(g3204), .b(n1112), .a(n1131) );
  nand2_812 NAND2_112 ( .c(I15993), .b(g10422), .a(I15992) );
  nand2_811 NAND2_113 ( .c(I5036), .b(g1019), .a(I5034) );
  nand2_810 NAND2_114 ( .c(I14263), .b(g8843), .a(g1814) );
  nand2_809 NAND2_115 ( .c(g8298), .b(I13249), .a(I13250) );
  nand2_808 NAND2_116 ( .c(I5135), .b(g521), .a(g525) );
  nand2_807 NAND2_117 ( .c(g2405), .b(I5485), .a(I5486) );
  nand2_806 NAND2_118 ( .c(I7034), .b(g3089), .a(I7033) );
  nand2_805 NAND2_119 ( .c(I15443), .b(g10007), .a(I15441) );
  nand2_804 NAND2_120 ( .c(I6166), .b(g2236), .a(g153) );
  nand2_803 NAND2_121 ( .c(I8624), .b(g4267), .a(g511) );
  nand2_802 NAND2_122 ( .c(I16015), .b(g10425), .a(n1339) );
  nand2_801 NAND2_123 ( .c(I8677), .b(g4374), .a(I8676) );
  nand2_800 NAND2_124 ( .c(I8576), .b(g4234), .a(I8575) );
  nand2_799 NAND2_125 ( .c(I14613), .b(g9204), .a(I14612) );
  nand2_798 NAND2_126 ( .c(I8716), .b(g4601), .a(I8715) );
  nand2_797 NAND2_127 ( .c(g3530), .b(I6715), .a(I6716) );
  nand2_796 NAND2_128 ( .c(g8405), .b(I13514), .a(I13515) );
  nand4_19 NAND4_2 ( .e(g4104), .d(g3215), .c(g3247), .b(g2439), .a(g3200) );
  nand2_795 NAND2_129 ( .c(I12003), .b(g5996), .a(I12002) );
  nand2_794 NAND2_130 ( .c(g2177), .b(I5127), .a(I5128) );
  nand2_793 NAND2_131 ( .c(g3010), .b(n1115), .a(n1130) );
  nand2_792 NAND2_132 ( .c(g5179), .b(I8576), .a(I8577) );
  nand2_791 NAND2_133 ( .c(I17395), .b(g11414), .a(I17393) );
  nand2_790 NAND2_134 ( .c(g7067), .b(I11279), .a(I11280) );
  nand4_18 NAND4_3 ( .e(g7994), .d(n1311), .c(g44), .b(n1309), .a(g42) );
  nand2_789 NAND2_135 ( .c(I6167), .b(g2236), .a(I6166) );
  nand2_788 NAND2_136 ( .c(I5265), .b(n1332), .a(I5263) );
  nand2_787 NAND2_137 ( .c(I6989), .b(g2760), .a(I6988) );
  nand2_786 NAND2_138 ( .c(I13274), .b(g8158), .a(I13272) );
  nand2_785 NAND2_139 ( .c(I10507), .b(g6221), .a(g786) );
  nand2_784 NAND2_140 ( .c(I13530), .b(g704), .a(I13529) );
  nand2_783 NAND2_141 ( .c(I5164), .b(g1508), .a(g1499) );
  nand2_782 NAND2_142 ( .c(g9107), .b(I14443), .a(I14444) );
  nand2_781 NAND2_143 ( .c(I9559), .b(g782), .a(I9557) );
  nand2_780 NAND2_144 ( .c(I8577), .b(g496), .a(I8575) );
  nand2_779 NAND2_145 ( .c(g2510), .b(I5592), .a(I5593) );
  nand2_778 NAND2_146 ( .c(g8177), .b(I13077), .a(I13078) );
  nand2_777 NAND2_147 ( .c(I8717), .b(g4052), .a(I8715) );
  nand2_776 NAND2_148 ( .c(I5296), .b(g794), .a(I5295) );
  nand2_775 NAND2_149 ( .c(g5209), .b(I8625), .a(I8626) );
  nand4_17 NAND4_4 ( .e(g7950), .d(g45), .c(g44), .b(g43), .a(n1308) );
  nand2_774 NAND2_150 ( .c(g2088), .b(I4911), .a(I4912) );
  nand2_773 NAND2_151 ( .c(I16000), .b(g10423), .a(I15999) );
  nand2_772 NAND2_152 ( .c(I5371), .b(g971), .a(g976) );
  nand2_771 NAND2_153 ( .c(g2215), .b(I5185), .a(I5186) );
  nand2_770 NAND2_154 ( .c(g7101), .b(n1270), .a(n1075) );
  nand2_769 NAND2_155 ( .c(I5675), .b(g1218), .a(g1223) );
  nand2_768 NAND2_156 ( .c(I8544), .b(g4218), .a(I8543) );
  nand2_767 NAND2_157 ( .c(g6577), .b(I10520), .a(I10521) );
  nand2_766 NAND2_158 ( .c(I5297), .b(g798), .a(I5295) );
  nand2_765 NAND2_159 ( .c(I13537), .b(g658), .a(g8157) );
  nand2_764 NAND2_160 ( .c(I13283), .b(g1927), .a(g8159) );
  nand2_763 NAND2_161 ( .c(g4749), .b(n1282), .a(n1131) );
  nand2_762 NAND2_162 ( .c(I11982), .b(g1482), .a(I11980) );
  nand2_761 NAND2_163 ( .c(I8514), .b(g4873), .a(I8513) );
  nand2_760 NAND2_164 ( .c(I13091), .b(g1840), .a(I13089) );
  nand2_759 NAND2_165 ( .c(g2943), .b(I6125), .a(I6126) );
  nand2_758 NAND2_166 ( .c(I15908), .b(g10302), .a(I15906) );
  nand2_757 NAND2_167 ( .c(I6879), .b(g3301), .a(g1351) );
  nand2_756 NAND2_168 ( .c(I8763), .b(g1129), .a(I8761) );
  nand2_755 NAND2_169 ( .c(I5449), .b(g1235), .a(g991) );
  nand3_21 NAND3_2 ( .d(g8825), .c(g8502), .b(g8738), .a(g8506) );
  nand2_754 NAND2_170 ( .c(I16007), .b(g10424), .a(g1776) );
  nand2_753 NAND2_171 ( .c(I5865), .b(g2107), .a(g2105) );
  nand2_752 NAND2_172 ( .c(I5604), .b(g1149), .a(g1153) );
  nand2_751 NAND2_173 ( .c(g2433), .b(I5517), .a(I5518) );
  nand2_750 NAND2_174 ( .c(I6111), .b(g1494), .a(I6109) );
  nand2_749 NAND2_175 ( .c(g2096), .b(I4929), .a(I4930) );
  nand2_748 NAND2_176 ( .c(I13522), .b(g695), .a(I13521) );
  nand2_747 NAND2_177 ( .c(I10770), .b(g5944), .a(I10769) );
  nand2_746 NAND2_178 ( .c(g6027), .b(n1269), .a(g4921) );
  nand4_16 NAND4_5 ( .e(g7992), .d(n1311), .c(g44), .b(n1309), .a(n1308) );
  nand2_745 NAND2_179 ( .c(I5539), .b(g1270), .a(I5538) );
  nand2_744 NAND2_180 ( .c(I17394), .b(g11415), .a(I17393) );
  nand2_743 NAND2_181 ( .c(I13553), .b(g668), .a(I13552) );
  nand2_742 NAND2_182 ( .c(I8642), .b(g516), .a(I8640) );
  nand2_741 NAND2_183 ( .c(g7573), .b(I12046), .a(I12047) );
  nand2_740 NAND2_184 ( .c(g11416), .b(I17296), .a(I17297) );
  nand2_739 NAND2_185 ( .c(g6003), .b(g5552), .a(g5548) );
  nand2_738 NAND2_186 ( .c(g8934), .b(I14278), .a(I14279) );
  nand2_737 NAND2_187 ( .c(I15992), .b(g10422), .a(n1333) );
  nand2_736 NAND2_188 ( .c(I7683), .b(g1023), .a(g3460) );
  nand2_735 NAND2_189 ( .c(I4910), .b(g386), .a(g318) );
  nand4_15 NAND4_6 ( .e(g3209), .d(n1149), .c(n1131), .b(n1109), .a(n1112) );
  nand2_734 NAND2_190 ( .c(I6794), .b(g143), .a(I6792) );
  nand2_733 NAND2_191 ( .c(I10521), .b(g822), .a(I10519) );
  nand2_732 NAND2_192 ( .c(I5486), .b(g1011), .a(I5484) );
  nand2_731 NAND2_193 ( .c(I15442), .b(g10013), .a(I15441) );
  nand2_730 NAND2_194 ( .c(g6858), .b(I10931), .a(I10932) );
  nand2_729 NAND2_195 ( .c(I5185), .b(g1415), .a(I5184) );
  nand2_728 NAND2_196 ( .c(g5304), .b(I8779), .a(I8780) );
  nand2_727 NAND2_197 ( .c(g2354), .b(g1515), .a(g1520) );
  nand2_726 NAND2_198 ( .c(I15615), .b(g10043), .a(g10153) );
  nand2_725 NAND2_199 ( .c(I17281), .b(g11221), .a(g11219) );
  nand2_724 NAND2_200 ( .c(I5470), .b(g999), .a(I5468) );
  nand2_723 NAND2_201 ( .c(I11509), .b(g6580), .a(I11508) );
  nand2_722 NAND2_202 ( .c(I5025), .b(g1275), .a(I5023) );
  nand2_721 NAND2_203 ( .c(I11508), .b(g6580), .a(g1806) );
  nand2_720 NAND2_204 ( .c(I15430), .b(g10001), .a(g9995) );
  nand2_719 NAND2_205 ( .c(I14612), .b(g9204), .a(g611) );
  nand2_718 NAND2_206 ( .c(g4675), .b(g4073), .a(g3247) );
  nand2_717 NAND2_207 ( .c(I14272), .b(g1822), .a(I14270) );
  nand2_716 NAND2_208 ( .c(g2979), .b(I6208), .a(I6209) );
  nand2_715 NAND2_209 ( .c(I17290), .b(g11223), .a(I17288) );
  nand2_714 NAND2_210 ( .c(g5269), .b(I8716), .a(I8717) );
  nand2_713 NAND2_211 ( .c(g4297), .b(I7563), .a(I7564) );
  nand2_712 NAND2_212 ( .c(I12002), .b(g5996), .a(g153) );
  nand2_711 NAND2_213 ( .c(I5006), .b(g421), .a(I5005) );
  nand2_710 NAND2_214 ( .c(I12128), .b(g170), .a(I12126) );
  nand2_709 NAND2_215 ( .c(I5105), .b(g431), .a(I5104) );
  nand2_708 NAND2_216 ( .c(I6323), .b(n1076), .a(I6322) );
  nand2_707 NAND2_217 ( .c(g7588), .b(I12093), .a(I12094) );
  nand2_706 NAND2_218 ( .c(I6666), .b(g2776), .a(I6664) );
  nand2_705 NAND2_219 ( .c(g3623), .b(I6761), .a(I6762) );
  nand2_704 NAND2_220 ( .c(I5373), .b(g976), .a(I5371) );
  nand2_703 NAND2_221 ( .c(I8529), .b(g481), .a(I8527) );
  nand2_702 NAND2_222 ( .c(I5283), .b(g758), .a(I5282) );
  nand2_701 NAND2_223 ( .c(I7224), .b(g2981), .a(I7223) );
  nand2_700 NAND2_224 ( .c(I5007), .b(g312), .a(I5005) );
  nand2_699 NAND2_225 ( .c(I5459), .b(g1240), .a(g1003) );
  nand2_698 NAND2_226 ( .c(I17297), .b(g11227), .a(I17295) );
  nand3_20 NAND3_3 ( .d(g8746), .c(g8289), .b(g47), .a(g46) );
  nand2_697 NAND2_227 ( .c(I6143), .b(n1157), .a(g646) );
  nand2_696 NAND2_228 ( .c(I5015), .b(g1011), .a(I5013) );
  nand2_695 NAND2_229 ( .c(g8932), .b(I14264), .a(I14265) );
  nand2_694 NAND2_230 ( .c(I16073), .b(g845), .a(I16072) );
  nand2_693 NAND2_231 ( .c(I6988), .b(g2760), .a(g986) );
  nand2_692 NAND2_232 ( .c(g3205), .b(g1814), .a(n1112) );
  nand2_691 NAND2_233 ( .c(I8652), .b(g778), .a(I8650) );
  nand2_690 NAND2_234 ( .c(I9558), .b(g5598), .a(I9557) );
  nand2_689 NAND2_235 ( .c(I5203), .b(g369), .a(I5202) );
  nand2_688 NAND2_236 ( .c(g7533), .b(I11936), .a(I11937) );
  nand2_687 NAND2_237 ( .c(g3634), .b(I6806), .a(I6807) );
  nand2_686 NAND2_238 ( .c(I6792), .b(g2959), .a(g143) );
  nand2_685 NAND2_239 ( .c(g3304), .b(I6468), .a(I6469) );
  nand2_684 NAND2_240 ( .c(I12145), .b(g158), .a(I12143) );
  nand2_683 NAND2_241 ( .c(g7596), .b(I12127), .a(I12128) );
  nand2_682 NAND2_242 ( .c(I13302), .b(g8162), .a(I13300) );
  nand2_681 NAND2_243 ( .c(I5502), .b(g1007), .a(I5500) );
  nand2_680 NAND2_244 ( .c(I9574), .b(g5608), .a(g818) );
  nand2_679 NAND2_245 ( .c(g3273), .b(I6448), .a(I6449) );
  nand2_678 NAND2_246 ( .c(I8670), .b(g4831), .a(I8669) );
  nand2_677 NAND2_247 ( .c(I7035), .b(g1868), .a(I7033) );
  nand2_676 NAND2_248 ( .c(I15453), .b(g10019), .a(I15451) );
  nand2_675 NAND2_249 ( .c(I8625), .b(g4267), .a(I8624) );
  nand2_674 NAND2_250 ( .c(I7876), .b(g4109), .a(I7875) );
  nand2_673 NAND2_251 ( .c(I14203), .b(g8825), .a(I14202) );
  nand2_672 NAND2_252 ( .c(I15607), .b(g10149), .a(g10144) );
  nand2_671 NAND2_253 ( .c(g2274), .b(I5324), .a(I5325) );
  nand2_670 NAND2_254 ( .c(I8740), .b(g1121), .a(I8738) );
  nand2_669 NAND2_255 ( .c(I17296), .b(g11229), .a(I17295) );
  nand2_668 NAND2_256 ( .c(g10507), .b(g10434), .a(g5859) );
  nand2_667 NAND2_257 ( .c(g2325), .b(g611), .a(g617) );
  nand2_666 NAND2_258 ( .c(I8606), .b(g506), .a(I8604) );
  nand2_665 NAND2_259 ( .c(I12087), .b(g1470), .a(I12085) );
  nand2_664 NAND2_260 ( .c(I13249), .b(g1891), .a(I13248) );
  nand2_663 NAND2_261 ( .c(I13248), .b(g1891), .a(g8148) );
  nand2_662 NAND2_262 ( .c(I13552), .b(g668), .a(g8262) );
  nand2_661 NAND2_263 ( .c(g2106), .b(I4979), .a(I4980) );
  nand2_660 NAND2_264 ( .c(I12069), .b(g139), .a(I12067) );
  nand2_659 NAND2_265 ( .c(g9204), .b(g6019), .a(g8942) );
  nand2_658 NAND2_266 ( .c(I12068), .b(g6045), .a(I12067) );
  nand2_657 NAND2_267 ( .c(I17503), .b(g11430), .a(g5269) );
  nand2_656 NAND2_268 ( .c(I7877), .b(g810), .a(I7875) );
  nand2_655 NAND2_269 ( .c(I5165), .b(g1508), .a(I5164) );
  nand2_654 NAND2_270 ( .c(g6740), .b(n1246), .a(n1149) );
  nand2_653 NAND2_271 ( .c(I6289), .b(g981), .a(I6287) );
  nand2_652 NAND2_272 ( .c(I6777), .b(g2892), .a(g650) );
  nand2_651 NAND2_273 ( .c(g5171), .b(I8562), .a(I8563) );
  nand2_650 NAND2_274 ( .c(I15891), .b(g853), .a(I15890) );
  nand2_649 NAND2_275 ( .c(I13090), .b(g8006), .a(I13089) );
  nand2_648 NAND2_276 ( .c(g11474), .b(I17460), .a(I17461) );
  nand4_14 NAND4_7 ( .e(g7942), .d(g45), .c(n1310), .b(g43), .a(g42) );
  nand2_647 NAND2_277 ( .c(I5538), .b(g1270), .a(g1023) );
  nand2_646 NAND2_278 ( .c(I7563), .b(g3533), .a(I7562) );
  nand2_645 NAND2_279 ( .c(I13513), .b(g686), .a(g8248) );
  nand2_644 NAND2_280 ( .c(g2107), .b(I4986), .a(I4987) );
  nand2_643 NAND2_281 ( .c(g2223), .b(I5203), .a(I5204) );
  nand2_642 NAND2_282 ( .c(I13505), .b(g677), .a(I13504) );
  nand2_641 NAND2_283 ( .c(I6209), .b(g802), .a(I6207) );
  nand2_640 NAND2_284 ( .c(I12086), .b(g5842), .a(I12085) );
  nand2_639 NAND2_285 ( .c(I8545), .b(g486), .a(I8543) );
  nand2_638 NAND2_286 ( .c(I8180), .b(g1786), .a(I8178) );
  nand2_637 NAND2_287 ( .c(g2115), .b(I5014), .a(I5015) );
  nand2_636 NAND2_288 ( .c(I8591), .b(g501), .a(I8589) );
  nand2_635 NAND2_289 ( .c(I10931), .b(g5863), .a(I10930) );
  nand2_634 NAND2_290 ( .c(I17402), .b(g11416), .a(I17400) );
  nand2_633 NAND2_291 ( .c(g8307), .b(I13294), .a(I13295) );
  nand2_632 NAND2_292 ( .c(I12144), .b(g6000), .a(I12143) );
  nand2_631 NAND2_293 ( .c(I10520), .b(g6231), .a(I10519) );
  nand2_630 NAND2_294 ( .c(I5263), .b(n1336), .a(n1332) );
  nand2_629 NAND2_295 ( .c(g8757), .b(n1241), .a(g4401) );
  nand2_628 NAND2_296 ( .c(I6714), .b(g2961), .a(g201) );
  nand2_627 NAND2_297 ( .c(I14211), .b(g599), .a(I14209) );
  nand2_626 NAND2_298 ( .c(I8515), .b(g3513), .a(I8513) );
  nand2_625 NAND2_299 ( .c(g2272), .b(I5316), .a(I5317) );
  nand2_624 NAND2_300 ( .c(I9946), .b(g5233), .a(g1796) );
  nand2_623 NAND2_301 ( .c(I8750), .b(g4613), .a(g1125) );
  nand2_622 NAND2_302 ( .c(I5605), .b(g1149), .a(I5604) );
  nand2_621 NAND2_303 ( .c(g8880), .b(I14203), .a(I14204) );
  nand2_620 NAND2_304 ( .c(I16051), .b(g837), .a(g10371) );
  nand2_619 NAND2_305 ( .c(I16072), .b(g845), .a(g10373) );
  nand2_618 NAND2_306 ( .c(g10440), .b(g10360), .a(g6037) );
  nand2_617 NAND2_307 ( .c(g8612), .b(I13858), .a(I13859) );
  nand2_616 NAND2_308 ( .c(I15872), .b(g1796), .a(I15870) );
  nand2_615 NAND2_309 ( .c(I8528), .b(g4879), .a(I8527) );
  nand2_614 NAND2_310 ( .c(g8629), .b(I13901), .a(I13902) );
  nand4_13 NAND4_8 ( .e(g8542), .d(n1112), .c(g1828), .b(g1814), .a(g8390) );
  nand2_613 NAND2_311 ( .c(I9947), .b(g5233), .a(I9946) );
  nand2_612 NAND2_312 ( .c(I6838), .b(g806), .a(I6836) );
  nand2_611 NAND2_313 ( .c(g7583), .b(I12068), .a(I12069) );
  nand2_610 NAND2_314 ( .c(g4803), .b(n1254), .a(n1386) );
  nand2_609 NAND2_315 ( .c(I17307), .b(g11231), .a(I17305) );
  nand2_608 NAND2_316 ( .c(g4538), .b(n1244), .a(n1130) );
  nand2_607 NAND2_317 ( .c(I15452), .b(g10025), .a(I15451) );
  nand2_606 NAND2_318 ( .c(I13857), .b(g8270), .a(g1448) );
  nand2_605 NAND2_319 ( .c(I14202), .b(g8825), .a(g591) );
  nand2_604 NAND2_320 ( .c(I13765), .b(g731), .a(g8417) );
  nand2_603 NAND2_321 ( .c(g2260), .b(I5296), .a(I5297) );
  nand4_12 NAND4_9 ( .e(g7986), .d(n1311), .c(n1310), .b(n1309), .a(g42) );
  nand2_602 NAND2_322 ( .c(g5226), .b(I8670), .a(I8671) );
  nand2_601 NAND2_323 ( .c(g8512), .b(n1279), .a(g8366) );
  nand2_600 NAND2_324 ( .c(I16046), .b(g10370), .a(I16044) );
  nand2_599 NAND2_325 ( .c(I13504), .b(g677), .a(g8247) );
  nand2_598 NAND2_326 ( .c(g10447), .b(g10363), .a(g5360) );
  nand2_597 NAND2_327 ( .c(g2167), .b(I5105), .a(I5106) );
  nand2_596 NAND2_328 ( .c(I8804), .b(g4677), .a(I8803) );
  nand2_595 NAND2_329 ( .c(g10472), .b(I16016), .a(I16017) );
  nand2_594 NAND2_330 ( .c(I17487), .b(g11474), .a(I17485) );
  nand2_593 NAND2_331 ( .c(I4995), .b(g416), .a(g309) );
  nand2_592 NAND2_332 ( .c(I12093), .b(g5810), .a(I12092) );
  nand4_11 NAND4_10 ( .e(g7987), .d(n1311), .c(n1310), .b(g43), .a(n1308) );
  nand2_591 NAND2_333 ( .c(g5227), .b(I8677), .a(I8678) );
  nand2_590 NAND2_334 ( .c(I5126), .b(g1386), .a(g1389) );
  nand2_589 NAND2_335 ( .c(g2321), .b(I5372), .a(I5373) );
  nand2_588 NAND2_336 ( .c(g7547), .b(I11974), .a(I11975) );
  nand2_587 NAND2_337 ( .c(I17306), .b(g11232), .a(I17305) );
  nand3_19 NAND3_4 ( .d(g6548), .c(g826), .b(g6124), .a(g6122) );
  nand2_586 NAND2_338 ( .c(I11995), .b(g6035), .a(g127) );
  nand2_585 NAND2_339 ( .c(I7225), .b(n1339), .a(I7223) );
  nand2_584 NAND2_340 ( .c(I11261), .b(g6775), .a(g826) );
  nand3_18 NAND3_5 ( .d(g8843), .c(g8542), .b(g8757), .a(g8545) );
  nand2_583 NAND2_341 ( .c(g2938), .b(I6110), .a(I6111) );
  nand2_582 NAND2_342 ( .c(I4942), .b(g396), .a(I4941) );
  nand2_581 NAND2_343 ( .c(g10394), .b(I15899), .a(I15900) );
  nand2_580 NAND2_344 ( .c(g8549), .b(g5527), .a(g8390) );
  nand2_579 NAND2_345 ( .c(g3070), .b(n1090), .a(g1206) );
  nand2_578 NAND2_346 ( .c(I4954), .b(g401), .a(g327) );
  nand2_577 NAND2_347 ( .c(I5023), .b(g995), .a(g1275) );
  nand2_576 NAND2_348 ( .c(g10446), .b(g10443), .a(g5350) );
  nand2_575 NAND2_349 ( .c(I16081), .b(g10374), .a(I16079) );
  nand2_574 NAND2_350 ( .c(I8641), .b(g4278), .a(I8640) );
  nand2_573 NAND2_351 ( .c(I6178), .b(g197), .a(I6176) );
  nand2_572 NAND2_352 ( .c(I12075), .b(g6015), .a(I12074) );
  nand2_571 NAND2_353 ( .c(I5127), .b(g1386), .a(I5126) );
  nand2_570 NAND2_354 ( .c(I5451), .b(g991), .a(I5449) );
  nand2_569 NAND2_355 ( .c(g4168), .b(I7322), .a(I7323) );
  nand2_568 NAND2_356 ( .c(I6288), .b(g2091), .a(I6287) );
  nand2_567 NAND2_357 ( .c(I8179), .b(g3685), .a(I8178) );
  nand2_566 NAND2_358 ( .c(I4912), .b(g318), .a(I4910) );
  nand2_565 NAND2_359 ( .c(I6805), .b(g3268), .a(n1334) );
  nand3_17 NAND3_6 ( .d(g3766), .c(g2439), .b(g3222), .a(g2493) );
  nand2_564 NAND2_360 ( .c(g3087), .b(I6288), .a(I6289) );
  nand2_563 NAND2_361 ( .c(I17486), .b(g11233), .a(I17485) );
  nand2_562 NAND2_362 ( .c(I4929), .b(g391), .a(I4928) );
  nand2_561 NAND2_363 ( .c(I15890), .b(g853), .a(g10286) );
  nand2_560 NAND2_364 ( .c(I16331), .b(n1201), .a(I16330) );
  nand2_559 NAND2_365 ( .c(I9575), .b(g5608), .a(I9574) );
  nand2_558 NAND2_366 ( .c(I13887), .b(g8267), .a(I13886) );
  nand2_557 NAND2_367 ( .c(g5308), .b(I8787), .a(I8788) );
  nand2_556 NAND2_368 ( .c(I13529), .b(g704), .a(g8253) );
  nand2_555 NAND2_369 ( .c(I6208), .b(g2534), .a(I6207) );
  nand2_554 NAND2_370 ( .c(g5217), .b(I8641), .a(I8642) );
  nand2_553 NAND2_371 ( .c(I5316), .b(g1032), .a(I5315) );
  nand2_552 NAND2_372 ( .c(g2111), .b(I5006), .a(I5007) );
  nand2_551 NAND2_373 ( .c(g10366), .b(g10285), .a(g5392) );
  nand2_550 NAND2_374 ( .c(I5034), .b(g1015), .a(g1019) );
  nand2_549 NAND2_375 ( .c(I13869), .b(g1403), .a(I13867) );
  nand2_548 NAND2_376 ( .c(I13868), .b(g8264), .a(I13867) );
  nand2_547 NAND2_377 ( .c(I15999), .b(g10423), .a(g1771) );
  nand2_546 NAND2_378 ( .c(I13259), .b(g1900), .a(I13258) );
  nand4_10 NAND4_11 ( .e(g3261), .d(n1155), .c(n1088), .b(n1078), .a(n1122) );
  nand2_545 NAND2_379 ( .c(g10481), .b(I16073), .a(I16074) );
  nand2_544 NAND2_380 ( .c(g2180), .b(I5136), .a(I5137) );
  nand3_16 NAND3_7 ( .d(g4976), .c(g2310), .b(g4604), .a(g3807) );
  nand2_543 NAND2_381 ( .c(g8506), .b(n1244), .a(g8366) );
  nand2_542 NAND2_382 ( .c(g2380), .b(I5460), .a(I5461) );
  nand2_541 NAND2_383 ( .c(I13258), .b(g1900), .a(g8153) );
  nand2_540 NAND2_384 ( .c(I5013), .b(g1007), .a(g1011) );
  nand2_539 NAND2_385 ( .c(g5196), .b(I8605), .a(I8606) );
  nand2_538 NAND2_386 ( .c(I10930), .b(g5863), .a(g5555) );
  nand2_537 NAND2_387 ( .c(I6770), .b(g3257), .a(g382) );
  nand2_536 NAND2_388 ( .c(g11449), .b(I17401), .a(I17402) );
  nand2_535 NAND2_389 ( .c(g11448), .b(I17394), .a(I17395) );
  nand2_534 NAND2_390 ( .c(I15717), .b(g10231), .a(I15716) );
  nand2_533 NAND2_391 ( .c(I5317), .b(g1027), .a(I5315) );
  nand2_532 NAND2_392 ( .c(I14210), .b(g8824), .a(I14209) );
  nand2_531 NAND2_393 ( .c(I17569), .b(g1610), .a(I17567) );
  nand2_530 NAND2_394 ( .c(I13878), .b(g1444), .a(I13876) );
  nand2_529 NAND2_395 ( .c(g8545), .b(n1282), .a(g8390) );
  nand2_528 NAND2_396 ( .c(g2515), .b(I5605), .a(I5606) );
  nand2_527 NAND2_397 ( .c(I14443), .b(g8970), .a(I14442) );
  nand2_526 NAND2_398 ( .c(g7557), .b(I11996), .a(I11997) );
  nand2_525 NAND2_399 ( .c(g8180), .b(I13090), .a(I13091) );
  nand2_524 NAND2_400 ( .c(I14279), .b(g1828), .a(I14277) );
  nand2_523 NAND2_401 ( .c(I17568), .b(g11496), .a(I17567) );
  nand2_522 NAND2_402 ( .c(I13886), .b(g8267), .a(g1440) );
  nand2_521 NAND2_403 ( .c(I7322), .b(g3047), .a(I7321) );
  nand2_520 NAND2_404 ( .c(I6990), .b(g986), .a(I6988) );
  nand2_519 NAND2_405 ( .c(I14278), .b(g8847), .a(I14277) );
  nand2_518 NAND2_406 ( .c(I7033), .b(g3089), .a(g1868) );
  nand2_517 NAND2_407 ( .c(I9006), .b(g4492), .a(g1791) );
  nand2_516 NAND2_408 ( .c(g8507), .b(n1280), .a(g8366) );
  nand2_515 NAND2_409 ( .c(I5460), .b(g1240), .a(I5459) );
  nand2_514 NAND2_410 ( .c(g4588), .b(n1264), .a(n1386) );
  nand2_513 NAND2_411 ( .c(I4986), .b(g999), .a(I4985) );
  nand3_15 NAND3_8 ( .d(g3247), .c(g1828), .b(n1109), .a(n1112) );
  nand2_512 NAND2_412 ( .c(I8651), .b(g4824), .a(I8650) );
  nand2_511 NAND2_413 ( .c(I13545), .b(g713), .a(I13544) );
  nand2_510 NAND2_414 ( .c(g8628), .b(I13894), .a(I13895) );
  nand2_509 NAND2_415 ( .c(I6138), .b(g378), .a(I6136) );
  nand2_508 NAND2_416 ( .c(I12074), .b(g6015), .a(g174) );
  nand2_507 NAND2_417 ( .c(g8630), .b(I13908), .a(I13909) );
  nand2_506 NAND2_418 ( .c(I13078), .b(g7963), .a(I13076) );
  nand2_505 NAND2_419 ( .c(I6109), .b(g2205), .a(g1494) );
  nand2_504 NAND2_420 ( .c(g8300), .b(I13259), .a(I13260) );
  nand2_503 NAND2_421 ( .c(I5501), .b(g1255), .a(I5500) );
  nand2_502 NAND2_422 ( .c(I17586), .b(n1293), .a(I17584) );
  nand2_501 NAND2_423 ( .c(I12092), .b(g5810), .a(g1490) );
  nand2_500 NAND2_424 ( .c(I13901), .b(g8261), .a(I13900) );
  nand2_499 NAND2_425 ( .c(I8795), .b(g4672), .a(g1145) );
  nand2_498 NAND2_426 ( .c(I6201), .b(g766), .a(I6199) );
  nand2_497 NAND2_427 ( .c(I14217), .b(g8826), .a(I14216) );
  nand2_496 NAND2_428 ( .c(I9007), .b(g4492), .a(I9006) );
  nand2_495 NAND2_429 ( .c(I13561), .b(g8263), .a(I13559) );
  nand2_494 NAND2_430 ( .c(I15716), .b(g10231), .a(g10229) );
  nand2_493 NAND2_431 ( .c(I6449), .b(g1776), .a(I6447) );
  nand2_492 NAND2_432 ( .c(I13295), .b(g8161), .a(I13293) );
  nand2_491 NAND2_433 ( .c(I4987), .b(g1003), .a(I4985) );
  nand2_490 NAND2_434 ( .c(I6715), .b(g2961), .a(I6714) );
  nand2_489 NAND2_435 ( .c(I17493), .b(g11430), .a(I17492) );
  nand2_488 NAND2_436 ( .c(I12215), .b(g7061), .a(I12214) );
  nand2_487 NAND2_437 ( .c(g2372), .b(I5450), .a(I5451) );
  nand2_486 NAND2_438 ( .c(g7062), .b(I11262), .a(I11263) );
  nand2_485 NAND2_439 ( .c(g2988), .b(I6225), .a(I6226) );
  nand2_484 NAND2_440 ( .c(I13309), .b(g617), .a(I13307) );
  nand2_483 NAND2_441 ( .c(g8839), .b(g8603), .a(g4401) );
  nand2_482 NAND2_442 ( .c(g2555), .b(I5676), .a(I5677) );
  nand2_481 NAND2_443 ( .c(g3662), .b(I6826), .a(I6827) );
  nand2_480 NAND2_444 ( .c(I13308), .b(g8190), .a(I13307) );
  nand2_479 NAND2_445 ( .c(g2792), .b(I5879), .a(I5880) );
  nand2_478 NAND2_446 ( .c(g4117), .b(g3041), .a(g3061) );
  nand2_477 NAND2_447 ( .c(I8543), .b(g4218), .a(g486) );
  nand2_476 NAND2_448 ( .c(g11549), .b(I17585), .a(I17586) );
  nand2_475 NAND2_449 ( .c(I6881), .b(g1351), .a(I6879) );
  nand2_474 NAND2_450 ( .c(I12138), .b(g131), .a(I12136) );
  nand2_473 NAND2_451 ( .c(I8729), .b(g4605), .a(I8728) );
  nand2_472 NAND2_452 ( .c(I14216), .b(g8826), .a(g605) );
  nand2_471 NAND2_453 ( .c(g10384), .b(I15871), .a(I15872) );
  nand2_470 NAND2_454 ( .c(I13260), .b(g8153), .a(I13258) );
  nand2_469 NAND2_455 ( .c(g2776), .b(I5866), .a(I5867) );
  nand2_468 NAND2_456 ( .c(I8513), .b(g4873), .a(g3513) );
  nand2_467 NAND2_457 ( .c(I13559), .b(g722), .a(g8263) );
  nand2_466 NAND2_458 ( .c(I8178), .b(g3685), .a(g1786) );
  nand2_465 NAND2_459 ( .c(g3631), .b(I6793), .a(I6794) );
  nand2_464 NAND2_460 ( .c(I6487), .b(g2306), .a(g1227) );
  nand2_463 NAND2_461 ( .c(I16080), .b(g849), .a(I16079) );
  nand2_462 NAND2_462 ( .c(I13893), .b(g8266), .a(g1436) );
  nand2_461 NAND2_463 ( .c(I12115), .b(g162), .a(I12113) );
  nand2_460 NAND2_464 ( .c(I6748), .b(g1453), .a(I6746) );
  nand2_459 NAND2_465 ( .c(I13544), .b(g713), .a(g8259) );
  nand2_458 NAND2_466 ( .c(I5484), .b(g1250), .a(g1011) );
  nand2_457 NAND2_467 ( .c(I4928), .b(g391), .a(g321) );
  nand2_456 NAND2_468 ( .c(I6226), .b(g1346), .a(I6224) );
  nand2_455 NAND2_469 ( .c(I8805), .b(g1113), .a(I8803) );
  nand2_454 NAND2_470 ( .c(I4930), .b(g321), .a(I4928) );
  nand2_453 NAND2_471 ( .c(I15880), .b(g1801), .a(I15878) );
  nand2_452 NAND2_472 ( .c(I14265), .b(g1814), .a(I14263) );
  nand2_451 NAND2_473 ( .c(I16031), .b(g829), .a(I16030) );
  nand2_450 NAND2_474 ( .c(g3585), .b(I6747), .a(I6748) );
  nand4_9 NAND4_12 ( .e(g3041), .d(n1075), .c(n1130), .b(n1126), .a(n1115) );
  nand2_449 NAND2_475 ( .c(g8933), .b(I14271), .a(I14272) );
  nand2_448 NAND2_476 ( .c(I16330), .b(n1201), .a(g4997) );
  nand2_447 NAND2_477 ( .c(I13267), .b(g8154), .a(I13265) );
  nand2_446 NAND2_478 ( .c(I13294), .b(g1882), .a(I13293) );
  nand2_445 NAND2_479 ( .c(g10231), .b(I15616), .a(I15617) );
  nand2_444 NAND2_480 ( .c(I14442), .b(g8970), .a(g1834) );
  nand2_443 NAND2_481 ( .c(I6793), .b(g2959), .a(I6792) );
  nand2_442 NAND2_482 ( .c(I4966), .b(g330), .a(I4964) );
  nand2_441 NAND2_483 ( .c(I8752), .b(g1125), .a(I8750) );
  nand2_440 NAND2_484 ( .c(I15432), .b(g9995), .a(I15430) );
  nand2_439 NAND2_485 ( .c(I12214), .b(g7061), .a(n1057) );
  nand2_438 NAND2_486 ( .c(g10511), .b(g10438), .a(g6032) );
  nand2_437 NAND2_487 ( .c(g3011), .b(g591), .a(n1115) );
  nand2_436 NAND2_488 ( .c(g5103), .b(I8480), .a(I8481) );
  nand2_435 NAND2_489 ( .c(I16087), .b(g861), .a(I16086) );
  nand2_434 NAND2_490 ( .c(g3734), .b(n1243), .a(g599) );
  nand2_433 NAND2_491 ( .c(I6664), .b(g2792), .a(g2776) );
  nand2_432 NAND2_492 ( .c(g8882), .b(I14217), .a(I14218) );
  nand2_431 NAND2_493 ( .c(I4955), .b(g401), .a(I4954) );
  nand2_430 NAND2_494 ( .c(I8786), .b(g4639), .a(g1141) );
  nand3_14 NAND3_9 ( .d(g3992), .c(n1112), .b(n1149), .a(g2990) );
  nand2_429 NAND2_495 ( .c(g10480), .b(I16066), .a(I16067) );
  nand2_428 NAND2_496 ( .c(I11915), .b(g5803), .a(I11914) );
  nand2_427 NAND2_497 ( .c(I8770), .b(g4619), .a(g1133) );
  nand2_426 NAND2_498 ( .c(I5516), .b(g1260), .a(g1019) );
  nand2_425 NAND2_499 ( .c(g8541), .b(n1291), .a(g8390) );
  nand2_424 NAND2_500 ( .c(I6188), .b(n1335), .a(I6186) );
  nand2_423 NAND2_501 ( .c(g5147), .b(I8544), .a(I8545) );
  nand3_13 NAND3_10 ( .d(g8744), .c(g8289), .b(g46), .a(n1313) );
  nand2_422 NAND2_502 ( .c(I5892), .b(g750), .a(I5891) );
  nand2_421 NAND2_503 ( .c(g8558), .b(I13766), .a(I13767) );
  nand2_420 NAND2_504 ( .c(I15258), .b(g9968), .a(I15256) );
  nand2_419 NAND2_505 ( .c(I13266), .b(g1909), .a(I13265) );
  nand2_418 NAND2_506 ( .c(I8787), .b(g4639), .a(I8786) );
  nand2_417 NAND2_507 ( .c(I6826), .b(g3281), .a(I6825) );
  nand2_416 NAND2_508 ( .c(I17283), .b(g11219), .a(I17281) );
  nand3_12 NAND3_11 ( .d(g5013), .c(g4749), .b(g3247), .a(g3205) );
  nand2_415 NAND2_509 ( .c(I17492), .b(g11430), .a(g3623) );
  nand2_414 NAND2_510 ( .c(g8511), .b(g5277), .a(g8366) );
  nand2_413 NAND2_511 ( .c(I16079), .b(g849), .a(g10374) );
  nand2_412 NAND2_512 ( .c(I5035), .b(g1015), .a(I5034) );
  nand2_411 NAND2_513 ( .c(I5517), .b(g1260), .a(I5516) );
  nand2_410 NAND2_514 ( .c(I7223), .b(g2981), .a(n1339) );
  nand2_409 NAND2_515 ( .c(I16086), .b(g861), .a(g10375) );
  nand2_408 NAND2_516 ( .c(g5317), .b(I8796), .a(I8797) );
  nand2_407 NAND2_517 ( .c(I15879), .b(g10359), .a(I15878) );
  nand2_406 NAND2_518 ( .c(I15878), .b(g10359), .a(g1801) );
  nand2_405 NAND2_519 ( .c(I12114), .b(g6002), .a(I12113) );
  nand2_404 NAND2_520 ( .c(I12107), .b(g6042), .a(I12106) );
  nand2_403 NAND2_521 ( .c(g2500), .b(g178), .a(g182) );
  nand2_402 NAND2_522 ( .c(I15994), .b(n1333), .a(I15992) );
  nand4_8 NAND4_13 ( .e(g7934), .d(g45), .c(n1310), .b(n1309), .a(g42) );
  nand2_401 NAND2_523 ( .c(g10469), .b(g10430), .a(g5999) );
  nand2_400 NAND2_524 ( .c(I14264), .b(g8843), .a(I14263) );
  nand2_399 NAND2_525 ( .c(I6448), .b(g2264), .a(I6447) );
  nand2_398 NAND2_526 ( .c(I13285), .b(g8159), .a(I13283) );
  nand2_397 NAND2_527 ( .c(g10468), .b(I16000), .a(I16001) );
  nand2_396 NAND2_528 ( .c(I6827), .b(g770), .a(I6825) );
  nand2_395 NAND2_529 ( .c(g8623), .b(I13877), .a(I13878) );
  nand2_394 NAND2_530 ( .c(I13900), .b(g8261), .a(g1428) );
  nand2_393 NAND2_531 ( .c(g2795), .b(I5892), .a(I5893) );
  nand2_392 NAND2_532 ( .c(I8575), .b(g4234), .a(g496) );
  nand2_391 NAND2_533 ( .c(I14209), .b(g8824), .a(g599) );
  nand2_390 NAND2_534 ( .c(I13560), .b(g722), .a(I13559) );
  nand2_389 NAND2_535 ( .c(I8715), .b(g4601), .a(g4052) );
  nand2_388 NAND2_536 ( .c(I8604), .b(g4259), .a(g506) );
  nand2_387 NAND2_537 ( .c(I16017), .b(n1339), .a(I16015) );
  nand2_386 NAND2_538 ( .c(I4941), .b(g396), .a(g324) );
  nand2_385 NAND2_539 ( .c(g2205), .b(I5165), .a(I5166) );
  nand3_11 NAND3_12 ( .d(g3753), .c(n1115), .b(n1075), .a(g2800) );
  nand2_384 NAND2_540 ( .c(I6467), .b(g23), .a(n1133) );
  nand2_383 NAND2_541 ( .c(I14614), .b(g611), .a(I14612) );
  nand2_382 NAND2_542 ( .c(g2104), .b(I4965), .a(I4966) );
  nand2_381 NAND2_543 ( .c(g2099), .b(I4942), .a(I4943) );
  nand2_380 NAND2_544 ( .c(I16023), .b(g10426), .a(g1786) );
  nand2_379 NAND2_545 ( .c(g10479), .b(I16059), .a(I16060) );
  nand3_10 NAND3_13 ( .d(g8737), .c(n1055), .b(g4921), .a(n1261) );
  nand2_378 NAND2_546 ( .c(g5942), .b(I9575), .a(I9576) );
  nand2_377 NAND2_547 ( .c(g10478), .b(I16052), .a(I16053) );
  nand2_376 NAND2_548 ( .c(I12004), .b(g153), .a(I12002) );
  nand2_375 NAND2_549 ( .c(I4911), .b(g386), .a(I4910) );
  nand2_374 NAND2_550 ( .c(I11914), .b(g5803), .a(g1494) );
  nand2_373 NAND2_551 ( .c(g7960), .b(g7409), .a(g5573) );
  nand2_372 NAND2_552 ( .c(I5295), .b(g794), .a(g798) );
  nand2_371 NAND2_553 ( .c(I12106), .b(g6042), .a(g135) );
  nand2_370 NAND2_554 ( .c(I8728), .b(g4605), .a(g1117) );
  nand2_369 NAND2_555 ( .c(g3681), .b(I6837), .a(I6838) );
  nand2_368 NAND2_556 ( .c(I11907), .b(g5838), .a(g1474) );
  nand2_367 NAND2_557 ( .c(I13907), .b(g8265), .a(g1432) );
  nand2_366 NAND2_558 ( .c(I8730), .b(g1117), .a(I8728) );
  nand2_365 NAND2_559 ( .c(g8551), .b(n1262), .a(g8390) );
  nand2_364 NAND2_560 ( .c(I4980), .b(g333), .a(I4978) );
  nand2_363 NAND2_561 ( .c(g2961), .b(I6177), .a(I6178) );
  nand2_362 NAND2_562 ( .c(g6019), .b(g617), .a(g4921) );
  nand2_361 NAND2_563 ( .c(I16016), .b(g10425), .a(I16015) );
  nand2_360 NAND2_564 ( .c(I11935), .b(g5857), .a(g1458) );
  nand2_359 NAND2_565 ( .c(I8678), .b(g1027), .a(I8676) );
  nand2_358 NAND2_566 ( .c(I17051), .b(g10923), .a(g11249) );
  nand2_357 NAND2_567 ( .c(g4482), .b(I7864), .a(I7865) );
  nand2_356 NAND2_568 ( .c(g7592), .b(I12107), .a(I12108) );
  nand2_355 NAND2_569 ( .c(g3460), .b(I6665), .a(I6666) );
  nand4_7 NAND4_14 ( .e(g7932), .d(g45), .c(n1310), .b(n1309), .a(n1308) );
  nand2_354 NAND2_570 ( .c(g7624), .b(I12215), .a(I12216) );
  nand4_6 NAND4_15 ( .e(g7953), .d(g45), .c(g44), .b(g43), .a(g42) );
  nand2_353 NAND2_571 ( .c(g8414), .b(I13553), .a(I13554) );
  nand2_352 NAND2_572 ( .c(I6168), .b(g153), .a(I6166) );
  nand2_351 NAND2_573 ( .c(I5229), .b(g182), .a(g148) );
  nand2_350 NAND2_574 ( .c(I6772), .b(g382), .a(I6770) );
  nand2_349 NAND2_575 ( .c(I16030), .b(g829), .a(g10368) );
  nand2_348 NAND2_576 ( .c(I13284), .b(g1927), .a(I13283) );
  nand2_347 NAND2_577 ( .c(I16065), .b(g10428), .a(g1806) );
  nand2_346 NAND2_578 ( .c(g2947), .b(I6137), .a(I6138) );
  nand2_345 NAND2_579 ( .c(I7321), .b(g3047), .a(g1231) );
  nand2_344 NAND2_580 ( .c(g2437), .b(I5529), .a(I5530) );
  nand2_343 NAND2_581 ( .c(g2102), .b(I4955), .a(I4956) );
  nand2_342 NAND2_582 ( .c(I17282), .b(g11221), .a(I17281) );
  nand2_341 NAND2_583 ( .c(I5620), .b(g1771), .a(I5618) );
  nand2_340 NAND2_584 ( .c(I8664), .b(g476), .a(I8662) );
  nand2_339 NAND2_585 ( .c(g7524), .b(I11915), .a(I11916) );
  nand2_338 NAND2_586 ( .c(g7717), .b(n1257), .a(g1950) );
  nand2_337 NAND2_587 ( .c(I16467), .b(g10716), .a(g10518) );
  nand2_336 NAND2_588 ( .c(I4972), .b(g991), .a(I4971) );
  nand2_335 NAND2_589 ( .c(I13554), .b(g8262), .a(I13552) );
  nand2_334 NAND2_590 ( .c(I16037), .b(g10427), .a(g1791) );
  nand2_333 NAND2_591 ( .c(g8302), .b(I13273), .a(I13274) );
  nand2_332 NAND2_592 ( .c(I4943), .b(g324), .a(I4941) );
  nand2_331 NAND2_593 ( .c(I5485), .b(g1250), .a(I5484) );
  nand2_330 NAND2_594 ( .c(g5527), .b(g3978), .a(g4749) );
  nand2_329 NAND2_595 ( .c(I10509), .b(g786), .a(I10507) );
  nand2_328 NAND2_596 ( .c(g7599), .b(I12144), .a(I12145) );
  nand2_327 NAND2_597 ( .c(I10508), .b(g6221), .a(I10507) );
  nand2_326 NAND2_598 ( .c(I6126), .b(g1419), .a(I6124) );
  nand2_325 NAND2_599 ( .c(I8671), .b(g814), .a(I8669) );
  nand2_324 NAND2_600 ( .c(I6760), .b(g2943), .a(g1448) );
  nand2_323 NAND2_601 ( .c(g3626), .b(I6778), .a(I6779) );
  nand2_322 NAND2_602 ( .c(I11973), .b(g5852), .a(g1462) );
  nand2_321 NAND2_603 ( .c(g2389), .b(I5469), .a(I5470) );
  nand2_320 NAND2_604 ( .c(I15617), .b(g10153), .a(I15615) );
  nand2_319 NAND2_605 ( .c(g5277), .b(g3734), .a(g4538) );
  nand2_318 NAND2_606 ( .c(I5005), .b(g421), .a(g312) );
  nand2_317 NAND2_607 ( .c(I6779), .b(g650), .a(I6777) );
  nand2_316 NAND2_608 ( .c(I6665), .b(g2792), .a(I6664) );
  nand2_315 NAND2_609 ( .c(I8589), .b(g4251), .a(g501) );
  nand2_314 NAND2_610 ( .c(g8412), .b(I13545), .a(I13546) );
  nand2_313 NAND2_611 ( .c(g2963), .b(I6187), .a(I6188) );
  nand2_312 NAND2_612 ( .c(I12045), .b(g5814), .a(g1486) );
  nand2_311 NAND2_613 ( .c(I16053), .b(g10371), .a(I16051) );
  nand2_310 NAND2_614 ( .c(g2109), .b(I4996), .a(I4997) );
  nand2_309 NAND2_615 ( .c(g11418), .b(I17306), .a(I17307) );
  nand2_308 NAND2_616 ( .c(I13539), .b(g8157), .a(I13537) );
  nand2_307 NAND2_617 ( .c(g10475), .b(I16031), .a(I16032) );
  nand2_306 NAND2_618 ( .c(I5324), .b(g1336), .a(I5323) );
  nand2_305 NAND2_619 ( .c(I13538), .b(g658), .a(I13537) );
  nand2_304 NAND2_620 ( .c(I5469), .b(g1245), .a(I5468) );
  nand2_303 NAND2_621 ( .c(I5540), .b(g1023), .a(I5538) );
  nand2_302 NAND2_622 ( .c(I17505), .b(g5269), .a(I17503) );
  nand2_301 NAND2_623 ( .c(I11241), .b(g6760), .a(g790) );
  nand2_300 NAND2_624 ( .c(I8803), .b(g4677), .a(g1113) );
  nand2_299 NAND2_625 ( .c(I12061), .b(g5824), .a(I12060) );
  nand2_298 NAND2_626 ( .c(I8780), .b(g1137), .a(I8778) );
  nand3_9 NAND3_14 ( .d(g8745), .c(g8289), .b(g47), .a(n1312) );
  nand2_297 NAND2_627 ( .c(I4979), .b(g411), .a(I4978) );
  nand2_296 NAND2_628 ( .c(g8109), .b(g48), .a(n1173) );
  nand2_295 NAND2_629 ( .c(g8309), .b(I13308), .a(I13309) );
  nand2_294 NAND2_630 ( .c(g6758), .b(I10770), .a(I10771) );
  nand2_293 NAND2_631 ( .c(I16009), .b(g1776), .a(I16007) );
  nand2_292 NAND2_632 ( .c(I15616), .b(g10043), .a(I15615) );
  nand2_291 NAND2_633 ( .c(I8662), .b(g4286), .a(g476) );
  nand2_290 NAND2_634 ( .c(I16008), .b(g10424), .a(I16007) );
  nand2_289 NAND2_635 ( .c(I13515), .b(g8248), .a(I13513) );
  nand2_288 NAND2_636 ( .c(I13991), .b(g622), .a(I13990) );
  nand2_287 NAND2_637 ( .c(g11276), .b(I17052), .a(I17053) );
  nand2_286 NAND2_638 ( .c(I15900), .b(g10287), .a(I15898) );
  nand2_285 NAND2_639 ( .c(g2419), .b(I5501), .a(I5502) );
  nand2_284 NAND2_640 ( .c(I16074), .b(g10373), .a(I16072) );
  nand2_283 NAND2_641 ( .c(I10769), .b(g5944), .a(g1801) );
  nand2_282 NAND2_642 ( .c(I7323), .b(g1231), .a(I7321) );
  nand2_281 NAND2_643 ( .c(g7978), .b(n1251), .a(g736) );
  nand2_280 NAND2_644 ( .c(I7875), .b(g4109), .a(g810) );
  nand2_279 NAND2_645 ( .c(I8562), .b(g4227), .a(I8561) );
  nand2_278 NAND2_646 ( .c(I15892), .b(g10286), .a(I15890) );
  nand2_277 NAND2_647 ( .c(g3771), .b(I6989), .a(I6990) );
  nand2_276 NAND2_648 ( .c(I8605), .b(g4259), .a(I8604) );
  nand2_275 NAND2_649 ( .c(g10153), .b(I15452), .a(I15453) );
  nand2_274 NAND2_650 ( .c(g5295), .b(I8762), .a(I8763) );
  nand2_273 NAND2_651 ( .c(I8751), .b(g4613), .a(I8750) );
  nand2_272 NAND2_652 ( .c(I15907), .b(g6899), .a(I15906) );
  nand2_271 NAND2_653 ( .c(I5136), .b(g521), .a(I5135) );
  nand2_270 NAND2_654 ( .c(I11263), .b(g826), .a(I11261) );
  nand2_269 NAND2_655 ( .c(I14204), .b(g591), .a(I14202) );
  nand2_268 NAND2_656 ( .c(g8881), .b(I14210), .a(I14211) );
  nand2_267 NAND2_657 ( .c(g2105), .b(I4972), .a(I4973) );
  nand3_8 NAND3_15 ( .d(g5557), .c(g4538), .b(g3071), .a(g3011) );
  nand2_266 NAND2_658 ( .c(I5230), .b(g182), .a(I5229) );
  nand2_265 NAND2_659 ( .c(I8669), .b(g4831), .a(g814) );
  nand2_264 NAND2_660 ( .c(g10474), .b(I16024), .a(I16025) );
  nand2_263 NAND2_661 ( .c(I8772), .b(g1133), .a(I8770) );
  nand2_262 NAND2_662 ( .c(g2445), .b(I5539), .a(I5540) );
  nand2_261 NAND2_663 ( .c(g8006), .b(g5552), .a(g7717) );
  nand2_260 NAND2_664 ( .c(I10932), .b(g5555), .a(I10930) );
  nand2_259 NAND2_665 ( .c(I17504), .b(g11430), .a(I17503) );
  nand2_258 NAND2_666 ( .c(I5137), .b(g525), .a(I5135) );
  nand2_257 NAND2_667 ( .c(g8305), .b(I13284), .a(I13285) );
  nand2_256 NAND2_668 ( .c(I5891), .b(g750), .a(n1144) );
  nand2_255 NAND2_669 ( .c(I13273), .b(g1918), .a(I13272) );
  nand2_254 NAND2_670 ( .c(I8480), .b(g4455), .a(I8479) );
  nand2_253 NAND2_671 ( .c(g4144), .b(g2160), .a(g109) );
  nand2_252 NAND2_672 ( .c(I15906), .b(g6899), .a(g10302) );
  nand2_251 NAND2_673 ( .c(I5342), .b(g315), .a(I5341) );
  nand2_250 NAND2_674 ( .c(I13514), .b(g686), .a(I13513) );
  nand2_249 NAND2_675 ( .c(g8407), .b(I13522), .a(I13523) );
  nand2_248 NAND2_676 ( .c(g4088), .b(I7224), .a(I7225) );
  nand2_247 NAND2_677 ( .c(g4488), .b(I7876), .a(I7877) );
  nand2_246 NAND2_678 ( .c(g7598), .b(I12137), .a(I12138) );
  nand3_7 NAND3_16 ( .d(g3222), .c(n1093), .b(g1814), .a(g1834) );
  nand2_245 NAND2_679 ( .c(I16052), .b(g837), .a(I16051) );
  nand2_244 NAND2_680 ( .c(I12127), .b(g6026), .a(I12126) );
  nand2_243 NAND2_681 ( .c(g10483), .b(I16087), .a(I16088) );
  nand2_242 NAND2_682 ( .c(g8415), .b(I13560), .a(I13561) );
  nand2_241 NAND2_683 ( .c(g11415), .b(I17289), .a(I17290) );
  nand2_240 NAND2_684 ( .c(g6573), .b(I10508), .a(I10509) );
  nand2_239 NAND2_685 ( .c(I5676), .b(g1218), .a(I5675) );
  nand2_238 NAND2_686 ( .c(I6778), .b(g2892), .a(I6777) );
  nand2_237 NAND2_687 ( .c(g9413), .b(I14613), .a(I14614) );
  nand2_236 NAND2_688 ( .c(I8779), .b(g4630), .a(I8778) );
  nand2_235 NAND2_689 ( .c(I5592), .b(g1696), .a(I5591) );
  nand4_5 NAND4_16 ( .e(g8502), .d(n1115), .c(g605), .b(g591), .a(g8366) );
  nand2_234 NAND2_690 ( .c(I15609), .b(g10144), .a(I15607) );
  nand2_233 NAND2_691 ( .c(I15608), .b(g10149), .a(I15607) );
  nand3_6 NAND3_17 ( .d(g3071), .c(g605), .b(n1126), .a(n1115) );
  nand2_232 NAND2_692 ( .c(g10509), .b(g10436), .a(g6023) );
  nand2_231 NAND2_693 ( .c(I17461), .b(g11448), .a(I17459) );
  nand2_230 NAND2_694 ( .c(I13506), .b(g8247), .a(I13504) );
  nand2_229 NAND2_695 ( .c(I5468), .b(g1245), .a(g999) );
  nand2_228 NAND2_696 ( .c(g5219), .b(I8651), .a(I8652) );
  nand2_227 NAND2_697 ( .c(I5677), .b(g1223), .a(I5675) );
  nand3_5 NAND3_18 ( .d(g8826), .c(g8512), .b(g8737), .a(g8648) );
  nand2_226 NAND2_698 ( .c(I17393), .b(g11415), .a(g11414) );
  nand2_225 NAND2_699 ( .c(I5866), .b(g2107), .a(I5865) );
  nand2_224 NAND2_700 ( .c(I12126), .b(g6026), .a(g170) );
  nand2_223 NAND2_701 ( .c(I4978), .b(g411), .a(g333) );
  nand2_222 NAND2_702 ( .c(g7587), .b(I12086), .a(I12087) );
  nand2_221 NAND2_703 ( .c(g5286), .b(I8751), .a(I8752) );
  nand2_220 NAND2_704 ( .c(g8308), .b(I13301), .a(I13302) );
  nand2_219 NAND2_705 ( .c(I7864), .b(g4099), .a(I7863) );
  nand2_218 NAND2_706 ( .c(I11981), .b(g5820), .a(I11980) );
  nand2_217 NAND2_707 ( .c(I12060), .b(g5824), .a(g1478) );
  nand2_216 NAND2_708 ( .c(g5225), .b(I8663), .a(I8664) );
  nand2_215 NAND2_709 ( .c(g11538), .b(I17568), .a(I17569) );
  nand2_214 NAND2_710 ( .c(I13767), .b(g8417), .a(I13765) );
  nand2_213 NAND2_711 ( .c(g10396), .b(I15907), .a(I15908) );
  nand2_212 NAND2_712 ( .c(I11262), .b(g6775), .a(I11261) );
  nand2_211 NAND2_713 ( .c(I13990), .b(g622), .a(n1261) );
  nand2_210 NAND2_714 ( .c(I6224), .b(g2544), .a(g1346) );
  nand2_209 NAND2_715 ( .c(I5867), .b(g2105), .a(I5865) );
  nand2_208 NAND2_716 ( .c(g2493), .b(g1834), .a(g1840) );
  nand2_207 NAND2_717 ( .c(I5893), .b(n1144), .a(I5891) );
  nand3_4 NAND3_19 ( .d(g3062), .c(n1099), .b(g591), .a(g611) );
  nand2_206 NAND2_718 ( .c(I13521), .b(g695), .a(g8249) );
  nand2_205 NAND2_719 ( .c(I5186), .b(g1515), .a(I5184) );
  nand2_204 NAND2_720 ( .c(I6771), .b(g3257), .a(I6770) );
  nand2_203 NAND2_721 ( .c(I5325), .b(g1341), .a(I5323) );
  nand2_202 NAND2_722 ( .c(I17459), .b(g11449), .a(g11448) );
  nand2_201 NAND2_723 ( .c(I9557), .b(g5598), .a(g782) );
  nand2_200 NAND2_724 ( .c(g11414), .b(I17282), .a(I17283) );
  nand2_199 NAND2_725 ( .c(I12067), .b(g6045), .a(g139) );
  nand2_198 NAND2_726 ( .c(I12094), .b(g1490), .a(I12092) );
  nand2_197 NAND2_727 ( .c(I4964), .b(g406), .a(g330) );
  nand2_196 NAND2_728 ( .c(I13272), .b(g1918), .a(g8158) );
  nand2_195 NAND2_729 ( .c(I9948), .b(g1796), .a(I9946) );
  nand2_194 NAND2_730 ( .c(g10302), .b(I15717), .a(I15718) );
  nand2_193 NAND2_731 ( .c(I16332), .b(g4997), .a(I16330) );
  nand2_192 NAND2_732 ( .c(I5106), .b(g435), .a(I5104) );
  nand2_191 NAND2_733 ( .c(g8847), .b(g8551), .a(g8683) );
  nand2_190 NAND2_734 ( .c(g2257), .b(I5283), .a(I5284) );
  nand2_189 NAND2_735 ( .c(I12019), .b(g6049), .a(g166) );
  nand2_188 NAND2_736 ( .c(I15441), .b(g10013), .a(g10007) );
  nand2_187 NAND2_737 ( .c(I11997), .b(g127), .a(I11995) );
  nand2_186 NAND2_738 ( .c(I8739), .b(g4607), .a(I8738) );
  nand2_185 NAND2_739 ( .c(I5461), .b(g1003), .a(I5459) );
  nand2_184 NAND2_740 ( .c(I13766), .b(g731), .a(I13765) );
  nand2_183 NAND2_741 ( .c(I8479), .b(g4455), .a(g3530) );
  nand2_182 NAND2_742 ( .c(I17295), .b(g11229), .a(g11227) );
  nand2_181 NAND2_743 ( .c(I14271), .b(g8840), .a(I14270) );
  nand2_180 NAND2_744 ( .c(I4971), .b(g991), .a(g995) );
  nand2_179 NAND2_745 ( .c(g8301), .b(I13266), .a(I13267) );
  nand2_178 NAND2_746 ( .c(I6110), .b(g2205), .a(I6109) );
  nand2_177 NAND2_747 ( .c(g10482), .b(I16080), .a(I16081) );
  nand2_176 NAND2_748 ( .c(g10779), .b(I16468), .a(I16469) );
  nand2_175 NAND2_749 ( .c(I6762), .b(g1448), .a(I6760) );
  nand2_174 NAND2_750 ( .c(I17289), .b(g11225), .a(I17288) );
  nand2_173 NAND2_751 ( .c(I5315), .b(g1032), .a(g1027) );
  nand2_172 NAND2_752 ( .c(I17288), .b(g11225), .a(g11223) );
  nand2_171 NAND2_753 ( .c(I13859), .b(g1448), .a(I13857) );
  nand2_170 NAND2_754 ( .c(g7548), .b(I11981), .a(I11982) );
  nand2_169 NAND2_755 ( .c(I13858), .b(g8270), .a(I13857) );
  nand2_168 NAND2_756 ( .c(I11996), .b(g6035), .a(I11995) );
  nand3_3 NAND3_20 ( .d(g8743), .c(g8289), .b(n1313), .a(n1312) );
  nand2_167 NAND2_757 ( .c(I5880), .b(g2115), .a(I5878) );
  nand2_166 NAND2_758 ( .c(g10513), .b(g10441), .a(g5345) );
  nand2_165 NAND2_759 ( .c(g8411), .b(I13538), .a(I13539) );
  nand2_164 NAND2_760 ( .c(I8626), .b(g511), .a(I8624) );
  nand2_163 NAND2_761 ( .c(g10505), .b(g10432), .a(g5938) );
  nand2_162 NAND2_762 ( .c(I5612), .b(g1280), .a(I5611) );
  nand2_161 NAND2_763 ( .c(g4821), .b(I8179), .a(I8180) );
  nand2_160 NAND2_764 ( .c(I12076), .b(g174), .a(I12074) );
  nand2_159 NAND2_765 ( .c(I12085), .b(g5842), .a(g1470) );
  nand2_158 NAND2_766 ( .c(g7567), .b(I12020), .a(I12021) );
  nand2_157 NAND2_767 ( .c(I5128), .b(g1389), .a(I5126) );
  nand2_156 NAND2_768 ( .c(I6489), .b(g1227), .a(I6487) );
  nand2_155 NAND2_769 ( .c(g7593), .b(I12114), .a(I12115) );
  nand2_154 NAND2_770 ( .c(I8778), .b(g4630), .a(g1137) );
  nand2_153 NAND2_771 ( .c(g10149), .b(I15442), .a(I15443) );
  nand2_152 NAND2_772 ( .c(I13902), .b(g1428), .a(I13900) );
  nand2_151 NAND2_773 ( .c(I13301), .b(g1936), .a(I13300) );
  nand2_150 NAND2_774 ( .c(g3215), .b(n1109), .a(g1822) );
  nand4_4 NAND4_17 ( .e(g7996), .d(n1311), .c(g44), .b(g43), .a(n1308) );
  nand2_149 NAND2_775 ( .c(I4985), .b(g999), .a(g1003) );
  nand2_148 NAND2_776 ( .c(I14444), .b(g1834), .a(I14442) );
  nand4_3 NAND4_18 ( .e(g8000), .d(n1311), .c(g44), .b(g43), .a(g42) );
  nand2_147 NAND2_777 ( .c(I5166), .b(g1499), .a(I5164) );
  nand2_146 NAND2_778 ( .c(I17460), .b(g11449), .a(I17459) );
  nand2_145 NAND2_779 ( .c(g3008), .b(n1066), .a(g878) );
  nand2_144 NAND2_780 ( .c(I6836), .b(g3287), .a(g806) );
  nand2_143 NAND2_781 ( .c(I5529), .b(g1265), .a(I5528) );
  nand2_142 NAND2_782 ( .c(g10229), .b(I15608), .a(I15609) );
  nand2_141 NAND2_783 ( .c(I13661), .b(g8322), .a(I13659) );
  nand2_140 NAND2_784 ( .c(I13895), .b(g1436), .a(I13893) );
  nand2_139 NAND2_785 ( .c(g2303), .b(I5342), .a(I5343) );
  nand2_138 NAND2_786 ( .c(I12039), .b(g5847), .a(I12038) );
  nand2_137 NAND2_787 ( .c(g5592), .b(I9007), .a(I9008) );
  nand2_136 NAND2_788 ( .c(I12038), .b(g5847), .a(g1466) );
  nand2_135 NAND2_789 ( .c(g3322), .b(I6488), .a(I6489) );
  nand2_134 NAND2_790 ( .c(I8561), .b(g4227), .a(g491) );
  nand2_133 NAND2_791 ( .c(I8527), .b(g4879), .a(g481) );
  nand2_132 NAND2_792 ( .c(I12143), .b(g6000), .a(g158) );
  nand2_131 NAND2_793 ( .c(I5619), .b(n1333), .a(I5618) );
  nand2_130 NAND2_794 ( .c(g10386), .b(I15879), .a(I15880) );
  nand2_129 NAND2_795 ( .c(I11980), .b(g5820), .a(g1482) );
  nand2_128 NAND2_796 ( .c(I6837), .b(g3287), .a(I6836) );
  nand2_127 NAND2_797 ( .c(I4973), .b(g995), .a(I4971) );
  nand2_126 NAND2_798 ( .c(I13888), .b(g1440), .a(I13886) );
  nand2_125 NAND2_799 ( .c(g7558), .b(I12003), .a(I12004) );
  nand2_124 NAND2_800 ( .c(I17494), .b(g3623), .a(I17492) );
  nand2_123 NAND2_801 ( .c(g11491), .b(I17493), .a(I17494) );
  nand2_122 NAND2_802 ( .c(I16045), .b(g833), .a(I16044) );
  nand2_121 NAND2_803 ( .c(I7684), .b(g1023), .a(I7683) );
  nand2_120 NAND2_804 ( .c(g4130), .b(g109), .a(n1057) );
  nand2_119 NAND2_805 ( .c(I8771), .b(g4619), .a(I8770) );
  nand2_118 NAND2_806 ( .c(I13546), .b(g8259), .a(I13544) );
  nand2_117 NAND2_807 ( .c(I13089), .b(g8006), .a(g1840) );
  nand2_116 NAND2_808 ( .c(g2117), .b(I5024), .a(I5025) );
  nand2_115 NAND2_809 ( .c(g5119), .b(I8514), .a(I8515) );
  nand2_114 NAND2_810 ( .c(g5319), .b(I8804), .a(I8805) );
  nand2_113 NAND2_811 ( .c(I15899), .b(g857), .a(I15898) );
  nand2_112 NAND2_812 ( .c(I5606), .b(g1153), .a(I5604) );
  nand2_111 NAND2_813 ( .c(I15898), .b(g857), .a(g10287) );
  nand2_110 NAND2_814 ( .c(I16032), .b(g10368), .a(I16030) );
  nand2_109 NAND2_815 ( .c(I17401), .b(g11418), .a(I17400) );
  nand2_108 NAND2_816 ( .c(I13659), .b(g1945), .a(g8322) );
  nand2_107 NAND2_817 ( .c(I8738), .b(g4607), .a(g1121) );
  nand2_106 NAND2_818 ( .c(I13250), .b(g8148), .a(I13248) );
  nand2_105 NAND2_819 ( .c(I15718), .b(g10229), .a(I15716) );
  nand2_104 NAND2_820 ( .c(I9008), .b(g1791), .a(I9006) );
  nand2_103 NAND2_821 ( .c(I6176), .b(g2177), .a(g197) );
  nand2_102 NAND2_822 ( .c(I7865), .b(g774), .a(I7863) );
  nand2_101 NAND2_823 ( .c(g5274), .b(I8729), .a(I8730) );
  nand2_100 NAND2_824 ( .c(I5341), .b(g315), .a(g426) );
  nand2_99 NAND2_825 ( .c(I17305), .b(g11232), .a(g11231) );
  nand2_98 NAND2_826 ( .c(I17053), .b(g11249), .a(I17051) );
  nand2_97 NAND2_827 ( .c(g5125), .b(I8528), .a(I8529) );
  nand2_96 NAND2_828 ( .c(I12216), .b(n1057), .a(I12214) );
  nand2_95 NAND2_829 ( .c(I6225), .b(g2544), .a(I6224) );
  nand2_94 NAND2_830 ( .c(I5879), .b(g2120), .a(I5878) );
  nand2_93 NAND2_831 ( .c(g3221), .b(g1834), .a(n1109) );
  nand2_92 NAND2_832 ( .c(I14270), .b(g8840), .a(g1822) );
  nand2_91 NAND2_833 ( .c(I6124), .b(g2215), .a(g1419) );
  nand2_90 NAND2_834 ( .c(I6324), .b(g1864), .a(I6322) );
  nand2_89 NAND2_835 ( .c(I13867), .b(g8264), .a(g1403) );
  nand2_88 NAND2_836 ( .c(I13894), .b(g8266), .a(I13893) );
  nand2_87 NAND2_837 ( .c(I6469), .b(n1133), .a(I6467) );
  nand2_86 NAND2_838 ( .c(I8663), .b(g4286), .a(I8662) );
  nand2_85 NAND2_839 ( .c(g7523), .b(I11908), .a(I11909) );
  nand2_84 NAND2_840 ( .c(I6177), .b(g2177), .a(I6176) );
  nand2_83 NAND2_841 ( .c(g5187), .b(I8590), .a(I8591) );
  nand2_82 NAND2_842 ( .c(I6287), .b(g2091), .a(g981) );
  nand2_81 NAND2_843 ( .c(I8762), .b(g4616), .a(I8761) );
  nand2_80 NAND2_844 ( .c(I15871), .b(g10358), .a(I15870) );
  nand3_2 NAND3_21 ( .d(g8840), .c(g8542), .b(g8541), .a(g8551) );
  nand2_79 NAND2_845 ( .c(g2250), .b(I5264), .a(I5265) );
  nand2_78 NAND2_846 ( .c(I8590), .b(g4251), .a(I8589) );
  nand2_77 NAND2_847 ( .c(I6199), .b(g2525), .a(g766) );
  nand2_76 NAND2_848 ( .c(I14218), .b(g605), .a(I14216) );
  nand2_75 NAND2_849 ( .c(g8190), .b(g6027), .a(g7978) );
  nand2_74 NAND2_850 ( .c(I5284), .b(g762), .a(I5282) );
  nand2_73 NAND2_851 ( .c(I17485), .b(g11233), .a(g11474) );
  nand2_72 NAND2_852 ( .c(I4965), .b(g406), .a(I4964) );
  nand2_71 NAND2_853 ( .c(I5591), .b(g1696), .a(g1703) );
  nand2_70 NAND2_854 ( .c(g8501), .b(n1292), .a(g8366) );
  nand2_69 NAND2_855 ( .c(I15451), .b(g10025), .a(g10019) );
  nand2_68 NAND2_856 ( .c(g8942), .b(g8823), .a(g4921) );
  nand2_67 NAND2_857 ( .c(I13877), .b(g8269), .a(I13876) );
  nand2_66 NAND2_858 ( .c(g7269), .b(I11509), .a(I11510) );
  nand2_65 NAND2_859 ( .c(I4996), .b(g416), .a(I4995) );
  nand2_64 NAND2_860 ( .c(I6144), .b(n1157), .a(I6143) );
  nand2_63 NAND2_861 ( .c(I17567), .b(g11496), .a(g1610) );
  nand2_62 NAND2_862 ( .c(g7572), .b(I12039), .a(I12040) );
  nand2_61 NAND2_863 ( .c(I6207), .b(g2534), .a(g802) );
  nand2_60 NAND2_864 ( .c(I14277), .b(g8847), .a(g1828) );
  nand2_59 NAND2_865 ( .c(I16059), .b(g841), .a(I16058) );
  nand2_58 NAND2_866 ( .c(I16025), .b(g1786), .a(I16023) );
  nand2_57 NAND2_867 ( .c(I8563), .b(g491), .a(I8561) );
  nand2_56 NAND2_868 ( .c(g3524), .b(g3209), .a(g3221) );
  nand2_55 NAND2_869 ( .c(I16058), .b(g841), .a(g10372) );
  nand2_54 NAND2_870 ( .c(I5204), .b(g374), .a(I5202) );
  nand2_53 NAND2_871 ( .c(I6488), .b(g2306), .a(I6487) );
  nand4_2 NAND4_19 ( .e(g3818), .d(g3056), .c(g3071), .b(g2310), .a(g3003) );
  nand2_52 NAND2_872 ( .c(I16044), .b(g833), .a(g10370) );
  nand2_51 NAND2_873 ( .c(g3717), .b(I6880), .a(I6881) );
  nand2_50 NAND2_874 ( .c(I13077), .b(g1872), .a(I13076) );
  nand2_49 NAND2_875 ( .c(g10043), .b(I15257), .a(I15258) );
  nand2_48 NAND2_876 ( .c(I11280), .b(g6485), .a(I11278) );
  nand2_47 NAND2_877 ( .c(I6825), .b(g3281), .a(g770) );
  nand2_46 NAND2_878 ( .c(I4997), .b(g309), .a(I4995) );
  nand2_45 NAND2_879 ( .c(I13300), .b(g1936), .a(g8162) );
  nand2_44 NAND2_880 ( .c(I5323), .b(g1336), .a(g1341) );
  nand2_43 NAND2_881 ( .c(I6136), .b(g2496), .a(g378) );
  nand2_42 NAND2_882 ( .c(g5935), .b(I9558), .a(I9559) );
  nand2_41 NAND2_883 ( .c(I5528), .b(g1265), .a(g1015) );
  nand2_40 NAND2_884 ( .c(I6806), .b(g3268), .a(I6805) );
  nand2_39 NAND2_885 ( .c(I5530), .b(g1015), .a(I5528) );
  nand2_38 NAND2_886 ( .c(g10886), .b(g10807), .a(g10805) );
  nand2_37 NAND2_887 ( .c(g3106), .b(I6323), .a(I6324) );
  nand2_36 NAND2_888 ( .c(I13876), .b(g8269), .a(g1444) );
  nand2_35 NAND2_889 ( .c(I6322), .b(n1076), .a(g1864) );
  nand2_34 NAND2_890 ( .c(g3061), .b(g611), .a(n1126) );
  nand2_33 NAND2_891 ( .c(g2439), .b(g1814), .a(g1828) );
  nand4_1 NAND4_20 ( .e(g7947), .d(g45), .c(g44), .b(n1309), .a(g42) );
  nand2_32 NAND2_892 ( .c(I9576), .b(g818), .a(I9574) );
  nand2_31 NAND2_893 ( .c(I13660), .b(g1945), .a(I13659) );
  nand2_30 NAND2_894 ( .c(g3200), .b(g1822), .a(n1131) );
  nand2_29 NAND2_895 ( .c(g4374), .b(I7684), .a(I7685) );
  nand2_28 NAND2_896 ( .c(I11916), .b(g1494), .a(I11914) );
  nand2_27 NAND2_897 ( .c(I5372), .b(g971), .a(I5371) );
  nand2_26 NAND2_898 ( .c(g3003), .b(g599), .a(n1130) );
  nand2_25 NAND2_899 ( .c(g8627), .b(I13887), .a(I13888) );
  nand2_24 NAND2_900 ( .c(I5618), .b(n1333), .a(g1771) );
  nand2_23 NAND2_901 ( .c(I6137), .b(g2496), .a(I6136) );
  nand2_22 NAND2_902 ( .c(I5343), .b(g426), .a(I5341) );
  nand2_21 NAND2_903 ( .c(I5282), .b(g758), .a(g762) );
  nand2_20 NAND2_904 ( .c(I13307), .b(g8190), .a(g617) );
  nand2_19 NAND2_905 ( .c(I13076), .b(g1872), .a(g7963) );
  nand2_18 NAND2_906 ( .c(I6807), .b(n1334), .a(I6805) );
  nand2_17 NAND2_907 ( .c(I11243), .b(g790), .a(I11241) );
  nand2_16 NAND2_908 ( .c(I17585), .b(g11217), .a(I17584) );
  nand2_15 NAND2_909 ( .c(I12137), .b(g6038), .a(I12136) );
  nand2_14 NAND2_910 ( .c(I7564), .b(g654), .a(I7562) );
  nand2_13 NAND2_911 ( .c(g2970), .b(I6200), .a(I6201) );
  nand2_12 NAND2_912 ( .c(g10144), .b(I15431), .a(I15432) );
  nand2_11 NAND2_913 ( .c(I8788), .b(g1141), .a(I8786) );
  nand2_10 NAND2_914 ( .c(g7054), .b(I11242), .a(I11243) );
  nand2_9 NAND2_915 ( .c(I17052), .b(g10923), .a(I17051) );
  nand2_8 NAND2_916 ( .c(g2120), .b(I5035), .a(I5036) );
  nand2_7 NAND2_917 ( .c(g8616), .b(I13868), .a(I13869) );
  nand2_6 NAND2_918 ( .c(I5202), .b(g369), .a(g374) );
  nand2_5 NAND2_919 ( .c(I16088), .b(g10375), .a(I16086) );
  nand2_4 NAND2_920 ( .c(I16024), .b(g10426), .a(I16023) );
  nand2_3 NAND2_921 ( .c(g11490), .b(I17486), .a(I17487) );
  nand2_2 NAND2_922 ( .c(I5518), .b(g1019), .a(I5516) );
  nand3_1 NAND3_22 ( .d(g5118), .c(g2439), .b(g4806), .a(g4073) );
  nand2_1 NAND2_923 ( .c(I12021), .b(g166), .a(I12019) );
  nor2_0 NOR2_0 ( .c(g6392), .b(g5859), .a(g5938) );
  nor2_97 NOR2_1 ( .c(g5938), .b(n1318), .a(n1392) );
  nor2_96 NOR2_2 ( .c(g2478), .b(g1610), .a(g1737) );
  nor2_95 NOR2_3 ( .c(g10374), .b(n1217), .a(n1392) );
  nor4_0 NOR4_0 ( .e(g4278), .d(n1079), .c(n1335), .b(n1332), .a(n1100) );
  nor2_94 NOR2_4 ( .c(g10424), .b(n1226), .a(n1392) );
  nor2_93 NOR2_5 ( .c(g10383), .b(n1226), .a(n1392) );
  nor2_92 NOR2_6 ( .c(g3118), .b(g2521), .a(g2514) );
  nor2_91 NOR2_7 ( .c(g9815), .b(n1321), .a(n1320) );
  nor2_90 NOR2_8 ( .c(g11077), .b(g10970), .a(g10971) );
  nor3_0 NOR3_0 ( .d(g9746), .c(n1327), .b(n1323), .a(n1331) );
  nor3_10 NOR3_1 ( .d(g3879), .c(n1160), .b(g2354), .a(g2353) );
  nor2_89 NOR2_9 ( .c(g10285), .b(n1218), .a(n1392) );
  nor2_88 NOR2_10 ( .c(g11480), .b(g11456), .a(n1164) );
  nor2_87 NOR2_11 ( .c(g4076), .b(g1707), .a(n1302) );
  nor2_86 NOR2_12 ( .c(g10570), .b(g10485), .a(g10324) );
  nor2_85 NOR2_13 ( .c(g10239), .b(g9317), .a(n1218) );
  nor2_84 NOR2_14 ( .c(g10594), .b(g10480), .a(g10521) );
  nor2_83 NOR2_15 ( .c(g9426), .b(g9052), .a(n1329) );
  nor2_82 NOR2_16 ( .c(g10382), .b(n1220), .a(n1392) );
  nor4_41 NOR4_1 ( .e(g4672), .d(n1104), .c(g1107), .b(g1104), .a(n1081) );
  nor2_81 NOR2_17 ( .c(g5360), .b(g105), .a(n1392) );
  nor4_40 NOR4_2 ( .e(g9387), .d(n1326), .c(n1330), .b(n1324), .a(I14596) );
  nor2_80 NOR2_18 ( .c(g10438), .b(n1219), .a(n1392) );
  nor4_39 NOR4_3 ( .e(g4613), .d(n1338), .c(n1141), .b(g1104), .a(g1101) );
  nor4_38 NOR4_4 ( .e(g9391), .d(n1326), .c(n1330), .b(n1324), .a(I14602) );
  nor3_9 NOR3_2 ( .d(g4572), .c(n1168), .b(n1181), .a(n1162) );
  nor3_8 NOR3_3 ( .d(g9757), .c(n1327), .b(n1323), .a(n1331) );
  nor2_79 NOR2_19 ( .c(g9416), .b(g9052), .a(n1329) );
  nor4_37 NOR4_5 ( .e(g9874), .d(g9519), .c(n1319), .b(g9579), .a(I15033) );
  nor2_78 NOR2_20 ( .c(g9654), .b(g9125), .a(n1328) );
  nor4_36 NOR4_6 ( .e(g9880), .d(g9751), .c(n1319), .b(g9557), .a(I15051) );
  nor4_35 NOR4_7 ( .e(g4873), .d(n1334), .c(n1335), .b(n1332), .a(n1100) );
  nor2_77 NOR2_21 ( .c(g2807), .b(n1386), .a(n1390) );
  nor2_76 NOR2_22 ( .c(g10441), .b(n1214), .a(n1392) );
  nor4_34 NOR4_8 ( .e(g4639), .d(n1104), .c(g1107), .b(g1104), .a(g1101) );
  nor2_75 NOR2_23 ( .c(g10435), .b(n1214), .a(n1392) );
  nor2_74 NOR2_24 ( .c(g10849), .b(g10739), .a(g2459) );
  nor4_33 NOR4_9 ( .e(g9606), .d(g9125), .c(g9111), .b(n1328), .a(n1325) );
  nor4_32 NOR4_10 ( .e(g9879), .d(g9747), .c(n1319), .b(g9566), .a(I15048) );
  nor2_73 NOR2_25 ( .c(g9506), .b(g9052), .a(n1329) );
  nor2_72 NOR2_26 ( .c(g6155), .b(g4974), .a(n1302) );
  nor2_71 NOR2_27 ( .c(g6355), .b(g6032), .a(g6023) );
  nor2_70 NOR2_28 ( .c(g9615), .b(g9052), .a(n1329) );
  nor2_69 NOR2_29 ( .c(g10371), .b(n1226), .a(n1392) );
  nor2_68 NOR2_30 ( .c(g9591), .b(g9125), .a(n1325) );
  nor2_67 NOR2_31 ( .c(g10359), .b(n1239), .a(n1392) );
  nor2_66 NOR2_32 ( .c(g10434), .b(n1226), .a(n1392) );
  nor2_65 NOR2_33 ( .c(g10358), .b(n1218), .a(n1392) );
  nor3_7 NOR3_4 ( .d(g9750), .c(n1327), .b(n1323), .a(n1331) );
  nor2_64 NOR2_34 ( .c(g10291), .b(n1218), .a(n1392) );
  nor4_31 NOR4_11 ( .e(g4227), .d(n1334), .c(n1098), .b(n1332), .a(n1336) );
  nor4_30 NOR4_12 ( .e(g9655), .d(n1326), .c(n1330), .b(n1324), .a(I14776) );
  nor4_29 NOR4_13 ( .e(g9410), .d(n1326), .c(n1330), .b(n1324), .a(I14607) );
  nor4_28 NOR4_14 ( .e(g9667), .d(g9125), .c(g9111), .b(n1328), .a(n1325) );
  nor2_63 NOR2_35 ( .c(g10563), .b(g10484), .a(g10322) );
  nor2_62 NOR2_36 ( .c(g9776), .b(n1321), .a(n1320) );
  nor2_61 NOR2_37 ( .c(g10324), .b(g9317), .a(n1217) );
  nor3_6 NOR3_5 ( .d(g4455), .c(n1183), .b(n1168), .a(n1181) );
  nor4_27 NOR4_15 ( .e(g9878), .d(g9754), .c(n1319), .b(g9560), .a(I15045) );
  nor2_60 NOR2_38 ( .c(g10360), .b(n1239), .a(n1392) );
  nor4_26 NOR4_16 ( .e(g9882), .d(g9742), .c(n1319), .b(g9563), .a(I15057) );
  nor2_59 NOR2_39 ( .c(g10370), .b(n1220), .a(n1392) );
  nor4_25 NOR4_17 ( .e(g4605), .d(n1338), .c(g1107), .b(n1052), .a(g1101) );
  nor2_58 NOR2_40 ( .c(g10420), .b(n1226), .a(n1392) );
  nor2_57 NOR2_41 ( .c(g10562), .b(g10483), .a(g10529) );
  nor2_56 NOR2_42 ( .c(g10427), .b(n1217), .a(n1392) );
  nor2_55 NOR2_43 ( .c(g5780), .b(n1062), .a(g4921) );
  nor2_54 NOR2_44 ( .c(g10385), .b(n1214), .a(n1392) );
  nor2_53 NOR2_45 ( .c(g10376), .b(n1217), .a(n1392) );
  nor2_52 NOR2_46 ( .c(g10426), .b(n1219), .a(n1392) );
  nor4_24 NOR4_18 ( .e(g4601), .d(n1338), .c(g1107), .b(g1104), .a(n1081) );
  nor2_51 NOR2_47 ( .c(g5573), .b(g4117), .a(g4432) );
  nor2_50 NOR2_48 ( .c(g9808), .b(n1321), .a(n1320) );
  nor2_49 NOR2_49 ( .c(g5999), .b(n1317), .a(n1392) );
  nor3_5 NOR3_6 ( .d(g9759), .c(n1327), .b(n1323), .a(n1331) );
  nor2_48 NOR2_50 ( .c(g6037), .b(n1101), .a(n1392) );
  nor2_47 NOR2_51 ( .c(g10287), .b(n1239), .a(n1392) );
  nor2_46 NOR2_52 ( .c(g5034), .b(g3524), .a(n1262) );
  nor4_23 NOR4_19 ( .e(g9362), .d(n1326), .c(n1330), .b(n1324), .a(I14585) );
  nor4_22 NOR4_20 ( .e(g9881), .d(g9516), .c(n1319), .b(g9573), .a(I15054) );
  nor2_45 NOR2_53 ( .c(g10443), .b(n1219), .a(n1392) );
  nor2_44 NOR2_54 ( .c(g10286), .b(n1218), .a(n1392) );
  nor3_4 NOR3_7 ( .d(g4276), .c(n1179), .b(g3261), .a(g2500) );
  nor4_21 NOR4_21 ( .e(g4616), .d(n1338), .c(n1141), .b(g1104), .a(n1081) );
  nor2_43 NOR2_55 ( .c(g10363), .b(n1217), .a(n1392) );
  nor2_42 NOR2_56 ( .c(g2862), .b(g2315), .a(g2305) );
  nor2_41 NOR2_57 ( .c(g10373), .b(n1219), .a(n1392) );
  nor2_40 NOR2_58 ( .c(g10423), .b(n1220), .a(n1392) );
  nor3_3 NOR3_8 ( .d(g9758), .c(n1327), .b(n1323), .a(n1331) );
  nor3_2 NOR3_9 ( .d(g9589), .c(g9125), .b(n1328), .a(n1325) );
  nor2_39 NOR2_59 ( .c(g9803), .b(n1321), .a(n1320) );
  nor2_38 NOR2_60 ( .c(g10430), .b(n1232), .a(n1392) );
  nor2_37 NOR2_61 ( .c(g9421), .b(g9052), .a(n1329) );
  nor2_36 NOR2_62 ( .c(g10362), .b(n1239), .a(n1392) );
  nor2_35 NOR2_63 ( .c(g2791), .b(n1114), .a(g750) );
  nor2_34 NOR2_64 ( .c(g9817), .b(n1321), .a(n1320) );
  nor4_20 NOR4_22 ( .e(g9605), .d(g9125), .c(g9111), .b(n1328), .a(n1325) );
  nor2_33 NOR2_65 ( .c(g10372), .b(n1214), .a(n1392) );
  nor2_32 NOR2_66 ( .c(g9669), .b(n1321), .a(n1320) );
  nor2_31 NOR2_67 ( .c(g10422), .b(n1232), .a(n1392) );
  nor2_30 NOR2_68 ( .c(g10436), .b(n1214), .a(n1392) );
  nor4_19 NOR4_23 ( .e(g5556), .d(n1189), .c(n1339), .b(n1064), .a(n1103) );
  nor4_18 NOR4_24 ( .e(g4286), .d(n1079), .c(n1335), .b(n1049), .a(n1336) );
  nor2_29 NOR2_69 ( .c(g4974), .b(g4502), .a(g3714) );
  nor2_28 NOR2_70 ( .c(g9779), .b(n1321), .a(n1320) );
  nor2_27 NOR2_71 ( .c(g9423), .b(g9052), .a(n1329) );
  nor2_26 NOR2_72 ( .c(g5350), .b(g3070), .a(n1392) );
  nor4_17 NOR4_25 ( .e(g9361), .d(n1326), .c(n1330), .b(n1324), .a(I14582) );
  nor4_16 NOR4_26 ( .e(g2459), .d(g1645), .c(g1642), .b(g1651), .a(g1648) );
  nor2_25 NOR2_73 ( .c(g10381), .b(n1232), .a(n1392) );
  nor4_15 NOR4_27 ( .e(g4259), .d(n1334), .c(n1098), .b(n1049), .a(n1100) );
  nor2_24 NOR2_74 ( .c(g10522), .b(g10401), .a(g10239) );
  nor2_23 NOR2_75 ( .c(g5392), .b(n1206), .a(n1392) );
  nor3_1 NOR3_10 ( .d(g4122), .c(n1204), .b(n1096), .a(g2538) );
  nor2_22 NOR2_76 ( .c(g6023), .b(n1054), .a(n1392) );
  nor2_21 NOR2_77 ( .c(g3462), .b(n1114), .a(g2795) );
  nor4_14 NOR4_28 ( .e(g4218), .d(n1334), .c(n1335), .b(n1049), .a(n1100) );
  nor4_13 NOR4_29 ( .e(g4267), .d(n1079), .c(n1335), .b(n1332), .a(n1336) );
  nor4_12 NOR4_30 ( .e(g4677), .d(n1104), .c(g1107), .b(n1052), .a(g1101) );
  nor2_20 NOR2_78 ( .c(g9646), .b(g9125), .a(n1325) );
  nor2_19 NOR2_79 ( .c(g2863), .b(g2316), .a(g2309) );
  nor4_11 NOR4_31 ( .e(g9616), .d(n1326), .c(n1330), .b(n1324), .a(I14751) );
  nor2_18 NOR2_80 ( .c(g6032), .b(g3008), .a(n1392) );
  nor4_10 NOR4_32 ( .e(g9647), .d(g9125), .c(g9111), .b(n1328), .a(n1325) );
  nor2_17 NOR2_81 ( .c(g5859), .b(g2987), .a(n1392) );
  nor2_16 NOR2_82 ( .c(g10433), .b(n1226), .a(n1392) );
  nor2_15 NOR2_83 ( .c(g10368), .b(n1232), .a(n1392) );
  nor4_9 NOR4_33 ( .e(g4251), .d(n1334), .c(n1098), .b(n1049), .a(n1336) );
  nor4_8 NOR4_34 ( .e(g9876), .d(g9522), .c(n1319), .b(g9052), .a(I15039) );
  nor4_7 NOR4_35 ( .e(g9656), .d(n1326), .c(n1330), .b(n1324), .a(I14779) );
  nor2_14 NOR2_84 ( .c(g8303), .b(g8209), .a(n1196) );
  nor2_13 NOR2_85 ( .c(g10429), .b(n1232), .a(n1392) );
  nor2_12 NOR2_86 ( .c(g10428), .b(n1232), .a(n1392) );
  nor4_6 NOR4_36 ( .e(g4234), .d(n1334), .c(n1098), .b(n1332), .a(n1100) );
  nor4_5 NOR4_37 ( .e(g9877), .d(g9512), .c(n1319), .b(g9569), .a(I15042) );
  nor2_11 NOR2_87 ( .c(g5186), .b(n1084), .a(g4401) );
  nor2_10 NOR2_88 ( .c(g9489), .b(g9052), .a(n1329) );
  nor4_4 NOR4_38 ( .e(g4619), .d(n1338), .c(n1141), .b(n1052), .a(g1101) );
  nor2_9 NOR2_89 ( .c(g10432), .b(n1220), .a(n1392) );
  nor2_8 NOR2_90 ( .c(g5345), .b(n1121), .a(n1392) );
  nor2_7 NOR2_91 ( .c(g5763), .b(g5350), .a(g5345) );
  nor2_6 NOR2_92 ( .c(g10375), .b(n1232), .a(n1392) );
  nor4_3 NOR4_39 ( .e(g4879), .d(n1334), .c(n1335), .b(n1049), .a(n1336) );
  nor4_2 NOR4_40 ( .e(g4607), .d(n1338), .c(g1107), .b(n1052), .a(n1081) );
  nor2_5 NOR2_93 ( .c(g10425), .b(n1214), .a(n1392) );
  nor2_4 NOR2_94 ( .c(g3107), .b(g2501), .a(g2499) );
  nor2_3 NOR2_95 ( .c(g10322), .b(g9317), .a(n1219) );
  nor4_1 NOR4_41 ( .e(g4630), .d(n1338), .c(n1141), .b(n1052), .a(n1081) );
  nor2_2 NOR2_96 ( .c(g10364), .b(n1220), .a(n1392) );
  nor2_1 NOR2_97 ( .c(g9781), .b(n1321), .a(n1320) );
  INVX1 U1097 ( .A(n1369), .Y(n1364) );
  INVX1 U1098 ( .A(n1368), .Y(n1366) );
  INVX1 U1099 ( .A(n1369), .Y(n1365) );
  INVX1 U1100 ( .A(n1374), .Y(n1363) );
  INVX1 U1101 ( .A(n1368), .Y(n1367) );
  INVX1 U1102 ( .A(g3015), .Y(n1368) );
  INVX1 U1103 ( .A(n1359), .Y(n1369) );
  INVX1 U1104 ( .A(n1360), .Y(n1382) );
  INVX1 U1105 ( .A(n1361), .Y(n1379) );
  INVX1 U1106 ( .A(n1360), .Y(n1377) );
  INVX1 U1107 ( .A(n1358), .Y(n1371) );
  INVX1 U1108 ( .A(n1360), .Y(n1378) );
  INVX1 U1109 ( .A(n1359), .Y(n1373) );
  INVX1 U1110 ( .A(n1359), .Y(n1375) );
  INVX1 U1111 ( .A(n1361), .Y(n1381) );
  INVX1 U1112 ( .A(n1358), .Y(n1372) );
  INVX1 U1113 ( .A(n1361), .Y(n1380) );
  INVX1 U1114 ( .A(n1359), .Y(n1374) );
  INVX1 U1115 ( .A(n1358), .Y(n1370) );
  INVX1 U1116 ( .A(n1360), .Y(n1376) );
  INVX1 U1117 ( .A(n1351), .Y(n1347) );
  INVX1 U1118 ( .A(n1350), .Y(n1348) );
  INVX1 U1119 ( .A(n1351), .Y(n1346) );
  INVX1 U1120 ( .A(n1350), .Y(n1349) );
  INVX1 U1121 ( .A(n1342), .Y(n1354) );
  INVX1 U1122 ( .A(n1343), .Y(n1353) );
  INVX1 U1123 ( .A(n1342), .Y(n1355) );
  INVX1 U1124 ( .A(n1343), .Y(n1356) );
  INVX1 U1125 ( .A(n1343), .Y(n1357) );
  INVX1 U1126 ( .A(g10950), .Y(n1177) );
  INVX1 U1127 ( .A(g11561), .Y(n1192) );
  INVX1 U1128 ( .A(g10809), .Y(n1163) );
  INVX1 U1129 ( .A(g8451), .Y(n1233) );
  INVX1 U1130 ( .A(g8488), .Y(n1213) );
  INVX1 U1131 ( .A(g7638), .Y(n1211) );
  INVX1 U1132 ( .A(g7246), .Y(n1210) );
  INVX1 U1133 ( .A(n1371), .Y(n1361) );
  INVX1 U1134 ( .A(n1362), .Y(n1359) );
  INVX1 U1135 ( .A(n1362), .Y(n1358) );
  INVX1 U1136 ( .A(n1373), .Y(n1360) );
  INVX1 U1137 ( .A(g10583), .Y(n1200) );
  INVX1 U1138 ( .A(g9331), .Y(n1190) );
  INVX1 U1139 ( .A(g9324), .Y(n1207) );
  BUFX3 U1140 ( .A(g9392), .Y(n1321) );
  BUFX3 U1141 ( .A(g9367), .Y(n1320) );
  INVX1 U1142 ( .A(n1341), .Y(n1350) );
  INVX1 U1143 ( .A(n1341), .Y(n1351) );
  INVX1 U1144 ( .A(n1344), .Y(n1342) );
  INVX1 U1145 ( .A(n1344), .Y(n1343) );
  INVX1 U1146 ( .A(n1341), .Y(n1352) );
  BUFX3 U1147 ( .A(g9536), .Y(n1319) );
  INVX1 U1148 ( .A(g10788), .Y(n1169) );
  INVX1 U1149 ( .A(g10937), .Y(n1191) );
  INVX1 U1150 ( .A(g10522), .Y(n1299) );
  INVX1 U1151 ( .A(n1327), .Y(n1182) );
  INVX1 U1152 ( .A(g10570), .Y(n1294) );
  INVX1 U1153 ( .A(g10385), .Y(n1297) );
  INVX1 U1154 ( .A(g8507), .Y(n1261) );
  INVX1 U1155 ( .A(g6488), .Y(n1245) );
  INVX1 U1156 ( .A(g8366), .Y(n1174) );
  INVX1 U1157 ( .A(g6740), .Y(n1257) );
  INVX1 U1158 ( .A(g7101), .Y(n1251) );
  INVX1 U1159 ( .A(g3041), .Y(n1264) );
  INVX1 U1160 ( .A(g3209), .Y(n1254) );
  INVX1 U1161 ( .A(g6003), .Y(n1253) );
  INVX1 U1162 ( .A(g2807), .Y(n1295) );
  INVX1 U1163 ( .A(g4977), .Y(n1180) );
  INVX1 U1164 ( .A(g5867), .Y(n1236) );
  INVX1 U1165 ( .A(g5309), .Y(n1216) );
  INVX1 U1166 ( .A(g3015), .Y(n1362) );
  INVX1 U1167 ( .A(g6351), .Y(n1173) );
  INVX1 U1168 ( .A(g9995), .Y(n1232) );
  INVX1 U1169 ( .A(g10013), .Y(n1214) );
  INVX1 U1170 ( .A(g10007), .Y(n1226) );
  INVX1 U1171 ( .A(g10019), .Y(n1219) );
  INVX1 U1172 ( .A(g10001), .Y(n1220) );
  INVX1 U1173 ( .A(g10025), .Y(n1217) );
  INVX1 U1174 ( .A(g9968), .Y(n1218) );
  INVX1 U1175 ( .A(g9974), .Y(n1239) );
  BUFX3 U1176 ( .A(g9240), .Y(n1330) );
  INVX1 U1177 ( .A(g8743), .Y(n1281) );
  BUFX3 U1178 ( .A(g9223), .Y(n1324) );
  BUFX3 U1179 ( .A(g9010), .Y(n1326) );
  INVX1 U1180 ( .A(g7947), .Y(n1290) );
  BUFX3 U1181 ( .A(g9173), .Y(n1328) );
  INVX1 U1182 ( .A(g11490), .Y(n1293) );
  INVX1 U1183 ( .A(n1345), .Y(n1341) );
  INVX1 U1184 ( .A(g10702), .Y(n1345) );
  INVX1 U1185 ( .A(g10702), .Y(n1344) );
  INVX1 U1186 ( .A(g7994), .Y(n1249) );
  INVX1 U1187 ( .A(g2303), .Y(n1285) );
  INVX1 U1188 ( .A(g3706), .Y(n1172) );
  BUFX3 U1189 ( .A(g9454), .Y(n1327) );
  INVX1 U1190 ( .A(g8746), .Y(n1255) );
  INVX1 U1191 ( .A(g11519), .Y(n1198) );
  INVX1 U1192 ( .A(g11276), .Y(n1275) );
  BUFX3 U1193 ( .A(g9151), .Y(n1325) );
  INVX1 U1194 ( .A(g9313), .Y(n1171) );
  BUFX3 U1195 ( .A(g9030), .Y(n1329) );
  INVX1 U1196 ( .A(g7950), .Y(n1250) );
  BUFX3 U1197 ( .A(g9292), .Y(n1331) );
  INVX1 U1198 ( .A(g7990), .Y(n1242) );
  BUFX3 U1199 ( .A(g9274), .Y(n1323) );
  INVX1 U1200 ( .A(g7987), .Y(n1260) );
  INVX1 U1201 ( .A(g2117), .Y(n1287) );
  INVX1 U1202 ( .A(g9052), .Y(n1340) );
  INVX1 U1203 ( .A(g7953), .Y(n1273) );
  INVX1 U1204 ( .A(g10563), .Y(n1296) );
  INVX1 U1205 ( .A(g10502), .Y(n1225) );
  INVX1 U1206 ( .A(g8546), .Y(n1241) );
  INVX1 U1207 ( .A(g3200), .Y(n1291) );
  INVX1 U1208 ( .A(g3003), .Y(n1292) );
  INVX1 U1209 ( .A(n1336), .Y(n1100) );
  INVX1 U1210 ( .A(g3753), .Y(n1269) );
  INVX1 U1211 ( .A(n1332), .Y(n1049) );
  INVX1 U1212 ( .A(n1335), .Y(n1098) );
  INVX1 U1213 ( .A(g8390), .Y(n1205) );
  INVX1 U1214 ( .A(n1334), .Y(n1079) );
  INVX1 U1215 ( .A(g3056), .Y(n1244) );
  INVX1 U1216 ( .A(g3374), .Y(n1164) );
  INVX1 U1217 ( .A(g3661), .Y(n1196) );
  INVX1 U1218 ( .A(g3101), .Y(n1183) );
  INVX1 U1219 ( .A(g5548), .Y(n1246) );
  INVX1 U1220 ( .A(g6019), .Y(n1270) );
  INVX1 U1221 ( .A(g3829), .Y(n1202) );
  INVX1 U1222 ( .A(g8574), .Y(n1224) );
  INVX1 U1223 ( .A(n1337), .Y(n1103) );
  INVX1 U1224 ( .A(g3992), .Y(n1265) );
  INVX1 U1225 ( .A(g5361), .Y(n1221) );
  INVX1 U1226 ( .A(g4640), .Y(n1229) );
  INVX1 U1227 ( .A(g4682), .Y(n1215) );
  INVX1 U1228 ( .A(n1322), .Y(n1199) );
  INVX1 U1229 ( .A(g3880), .Y(n1159) );
  INVX1 U1230 ( .A(g5557), .Y(n1276) );
  INVX1 U1231 ( .A(g5013), .Y(n1267) );
  INVX1 U1232 ( .A(n1338), .Y(n1104) );
  INVX1 U1233 ( .A(g3247), .Y(n1262) );
  INVX1 U1234 ( .A(n1388), .Y(n1386) );
  INVX1 U1235 ( .A(g5405), .Y(n1231) );
  INVX1 U1236 ( .A(g5576), .Y(n1234) );
  INVX1 U1237 ( .A(g9257), .Y(n1197) );
  INVX1 U1238 ( .A(g9268), .Y(n1186) );
  INVX1 U1239 ( .A(g9271), .Y(n1175) );
  INVX1 U1240 ( .A(g9256), .Y(n1195) );
  INVX1 U1241 ( .A(g3215), .Y(n1282) );
  INVX1 U1242 ( .A(g3071), .Y(n1279) );
  INVX1 U1243 ( .A(g2459), .Y(n1298) );
  INVX1 U1244 ( .A(g4117), .Y(n1263) );
  INVX1 U1245 ( .A(g3524), .Y(n1288) );
  INVX1 U1246 ( .A(g3062), .Y(n1280) );
  INVX1 U1247 ( .A(g3222), .Y(n1278) );
  INVX1 U1248 ( .A(g3108), .Y(n1181) );
  INVX1 U1249 ( .A(n1389), .Y(g2355) );
  INVX1 U1250 ( .A(g3104), .Y(n1168) );
  INVX1 U1251 ( .A(g8289), .Y(n1184) );
  INVX1 U1252 ( .A(g3120), .Y(n1228) );
  INVX1 U1253 ( .A(g2744), .Y(n1222) );
  INVX1 U1254 ( .A(g7624), .Y(n1272) );
  INVX1 U1255 ( .A(g4421), .Y(n1176) );
  INVX1 U1256 ( .A(g3111), .Y(n1162) );
  INVX1 U1257 ( .A(g3586), .Y(n1161) );
  INVX1 U1258 ( .A(g2276), .Y(n1206) );
  INVX1 U1259 ( .A(g4144), .Y(n1277) );
  INVX1 U1260 ( .A(g3863), .Y(n1185) );
  INVX1 U1261 ( .A(g7671), .Y(n1247) );
  INVX1 U1262 ( .A(g4089), .Y(n1227) );
  INVX1 U1263 ( .A(n1333), .Y(n1067) );
  INVX1 U1264 ( .A(n1384), .Y(n1383) );
  INVX1 U1265 ( .A(g7942), .Y(n1258) );
  INVX1 U1266 ( .A(g30), .Y(n1305) );
  INVX1 U1267 ( .A(g8745), .Y(n1274) );
  INVX1 U1268 ( .A(g8744), .Y(n1266) );
  INVX1 U1269 ( .A(g11580), .Y(n1212) );
  INVX1 U1270 ( .A(g48), .Y(n1385) );
  INVX1 U1271 ( .A(g41), .Y(n1307) );
  INVX1 U1272 ( .A(g45), .Y(n1311) );
  INVX1 U1273 ( .A(g7992), .Y(n1252) );
  INVX1 U1274 ( .A(g43), .Y(n1309) );
  INVX1 U1275 ( .A(g44), .Y(n1310) );
  INVX1 U1276 ( .A(g42), .Y(n1308) );
  INVX1 U1277 ( .A(g7996), .Y(n1283) );
  INVX1 U1278 ( .A(g7932), .Y(n1271) );
  INVX1 U1279 ( .A(g8000), .Y(n1284) );
  INVX1 U1280 ( .A(g7934), .Y(n1268) );
  INVX1 U1281 ( .A(g47), .Y(n1313) );
  INVX1 U1282 ( .A(g46), .Y(n1312) );
  INVX1 U1283 ( .A(g31), .Y(n1306) );
  INVX1 U1284 ( .A(g10334), .Y(n1194) );
  INVX1 U1285 ( .A(g10268), .Y(n1187) );
  INVX1 U1286 ( .A(g10740), .Y(n1193) );
  INVX1 U1287 ( .A(g10357), .Y(n1201) );
  INVX1 U1288 ( .A(g1811), .Y(n1142) );
  INVX1 U1289 ( .A(g10331), .Y(n1203) );
  INVX1 U1290 ( .A(g1854), .Y(n1116) );
  INVX1 U1291 ( .A(g10328), .Y(n1167) );
  INVX1 U1292 ( .A(g10325), .Y(n1170) );
  INVX1 U1293 ( .A(g10348), .Y(n1165) );
  INVX1 U1294 ( .A(g10333), .Y(n1166) );
  INVX1 U1295 ( .A(g654), .Y(n1091) );
  INVX1 U1296 ( .A(g599), .Y(n1115) );
  INVX1 U1297 ( .A(g591), .Y(n1126) );
  INVX1 U1298 ( .A(g650), .Y(n1140) );
  INVX1 U1299 ( .A(g646), .Y(n1059) );
  INVX1 U1300 ( .A(g7067), .Y(n1248) );
  BUFX3 U1301 ( .A(g471), .Y(n1334) );
  INVX1 U1302 ( .A(g2310), .Y(n1243) );
  INVX1 U1303 ( .A(g109), .Y(n1392) );
  BUFX3 U1304 ( .A(g466), .Y(n1335) );
  BUFX3 U1305 ( .A(g456), .Y(n1336) );
  BUFX3 U1306 ( .A(g461), .Y(n1332) );
  INVX1 U1307 ( .A(g643), .Y(n1157) );
  INVX1 U1308 ( .A(g1900), .Y(n1120) );
  INVX1 U1309 ( .A(g686), .Y(n1117) );
  INVX1 U1310 ( .A(g1909), .Y(n1150) );
  INVX1 U1311 ( .A(g695), .Y(n1048) );
  INVX1 U1312 ( .A(g1918), .Y(n1111) );
  INVX1 U1313 ( .A(g704), .Y(n1058) );
  INVX1 U1314 ( .A(g1927), .Y(n1056) );
  INVX1 U1315 ( .A(g713), .Y(n1047) );
  INVX1 U1316 ( .A(g1936), .Y(n1092) );
  INVX1 U1317 ( .A(g722), .Y(n1106) );
  INVX1 U1318 ( .A(g1891), .Y(n1125) );
  INVX1 U1319 ( .A(g677), .Y(n1148) );
  INVX1 U1320 ( .A(g1882), .Y(n1045) );
  INVX1 U1321 ( .A(g668), .Y(n1135) );
  INVX1 U1322 ( .A(g7986), .Y(n1259) );
  INVX1 U1323 ( .A(g1872), .Y(n1147) );
  INVX1 U1324 ( .A(g658), .Y(n1137) );
  INVX1 U1325 ( .A(g731), .Y(n1127) );
  INVX1 U1326 ( .A(g1945), .Y(n1102) );
  INVX1 U1327 ( .A(g1868), .Y(n1069) );
  INVX1 U1328 ( .A(g1357), .Y(n1097) );
  INVX1 U1329 ( .A(g876), .Y(n1066) );
  INVX1 U1330 ( .A(g1101), .Y(n1081) );
  INVX1 U1331 ( .A(g1104), .Y(n1052) );
  INVX1 U1332 ( .A(g1822), .Y(n1112) );
  INVX1 U1333 ( .A(g1107), .Y(n1141) );
  INVX1 U1334 ( .A(g2563), .Y(n1160) );
  INVX1 U1335 ( .A(g1453), .Y(n1096) );
  INVX1 U1336 ( .A(g2161), .Y(n1204) );
  INVX1 U1337 ( .A(g1718), .Y(n1071) );
  INVX1 U1338 ( .A(g1814), .Y(n1109) );
  INVX1 U1339 ( .A(g605), .Y(n1130) );
  INVX1 U1340 ( .A(g1828), .Y(n1131) );
  INVX1 U1341 ( .A(g1864), .Y(n1050) );
  BUFX3 U1342 ( .A(g4807), .Y(n1322) );
  INVX1 U1343 ( .A(g1713), .Y(n1083) );
  INVX1 U1344 ( .A(g2439), .Y(n1289) );
  INVX1 U1345 ( .A(g611), .Y(n1075) );
  INVX1 U1346 ( .A(g1834), .Y(n1149) );
  INVX1 U1347 ( .A(g127), .Y(n1156) );
  INVX1 U1348 ( .A(g1861), .Y(n1076) );
  BUFX3 U1349 ( .A(g1110), .Y(n1338) );
  BUFX3 U1350 ( .A(g1690), .Y(n1337) );
  BUFX3 U1351 ( .A(g1766), .Y(n1333) );
  INVX1 U1352 ( .A(g153), .Y(n1078) );
  INVX1 U1353 ( .A(g1840), .Y(n1093) );
  INVX1 U1354 ( .A(g617), .Y(n1099) );
  INVX1 U1355 ( .A(g622), .Y(n1055) );
  BUFX3 U1356 ( .A(g1781), .Y(n1339) );
  INVX1 U1357 ( .A(g639), .Y(n1062) );
  INVX1 U1358 ( .A(g1857), .Y(n1084) );
  INVX1 U1359 ( .A(g148), .Y(n1122) );
  INVX1 U1360 ( .A(g201), .Y(n1139) );
  INVX1 U1361 ( .A(g1389), .Y(n1060) );
  INVX1 U1362 ( .A(g197), .Y(n1143) );
  INVX1 U1363 ( .A(g636), .Y(n1128) );
  INVX1 U1364 ( .A(g1703), .Y(n1132) );
  INVX1 U1365 ( .A(g12), .Y(n1158) );
  INVX1 U1366 ( .A(g143), .Y(n1108) );
  INVX1 U1367 ( .A(g192), .Y(n1105) );
  INVX1 U1368 ( .A(g248), .Y(n1063) );
  INVX1 U1369 ( .A(g131), .Y(n1146) );
  INVX1 U1370 ( .A(g18), .Y(n1390) );
  INVX1 U1371 ( .A(g18), .Y(n1389) );
  INVX1 U1372 ( .A(g18), .Y(n1391) );
  INVX1 U1373 ( .A(g139), .Y(n1136) );
  INVX1 U1374 ( .A(g18), .Y(n1388) );
  INVX1 U1375 ( .A(g135), .Y(n1152) );
  INVX1 U1376 ( .A(g2794), .Y(n1179) );
  INVX1 U1377 ( .A(g1374), .Y(n1153) );
  INVX1 U1378 ( .A(g115), .Y(n1151) );
  INVX1 U1379 ( .A(g119), .Y(n1134) );
  INVX1 U1380 ( .A(g231), .Y(n1086) );
  INVX1 U1381 ( .A(g219), .Y(n1073) );
  INVX1 U1382 ( .A(g225), .Y(n1074) );
  INVX1 U1383 ( .A(g237), .Y(n1113) );
  INVX1 U1384 ( .A(g243), .Y(n1053) );
  INVX1 U1385 ( .A(g1696), .Y(n1301) );
  INVX1 U1386 ( .A(g1368), .Y(n1082) );
  INVX1 U1387 ( .A(g1362), .Y(n1065) );
  INVX1 U1388 ( .A(g1361), .Y(n1090) );
  INVX1 U1389 ( .A(g882), .Y(n1072) );
  INVX1 U1390 ( .A(g3423), .Y(n1189) );
  INVX1 U1391 ( .A(g757), .Y(n1054) );
  INVX1 U1392 ( .A(g108), .Y(n1121) );
  INVX1 U1393 ( .A(g881), .Y(n1318) );
  INVX1 U1394 ( .A(g85), .Y(n1316) );
  INVX1 U1395 ( .A(g3304), .Y(n1256) );
  INVX1 U1396 ( .A(g4130), .Y(n1286) );
  INVX1 U1397 ( .A(g590), .Y(n1057) );
  INVX1 U1398 ( .A(g754), .Y(n1144) );
  INVX1 U1399 ( .A(g746), .Y(n1114) );
  INVX1 U1400 ( .A(g1700), .Y(n1302) );
  INVX1 U1401 ( .A(g627), .Y(n1089) );
  INVX1 U1402 ( .A(g26), .Y(n1133) );
  INVX1 U1403 ( .A(g1707), .Y(n1064) );
  INVX1 U1404 ( .A(g3688), .Y(n1223) );
  INVX1 U1405 ( .A(g7651), .Y(n1237) );
  INVX1 U1406 ( .A(g7664), .Y(n1209) );
  INVX1 U1407 ( .A(g114), .Y(n1145) );
  INVX1 U1408 ( .A(g3354), .Y(n1235) );
  INVX1 U1409 ( .A(g4300), .Y(n1240) );
  INVX1 U1410 ( .A(g3698), .Y(n1208) );
  INVX1 U1411 ( .A(g7712), .Y(n1238) );
  INVX1 U1412 ( .A(g158), .Y(n1088) );
  INVX1 U1413 ( .A(g162), .Y(n1155) );
  INVX1 U1414 ( .A(g1845), .Y(n1124) );
  INVX1 U1415 ( .A(g794), .Y(n1094) );
  INVX1 U1416 ( .A(g1212), .Y(n1110) );
  INVX1 U1417 ( .A(g971), .Y(n1107) );
  INVX1 U1418 ( .A(g1336), .Y(n1123) );
  INVX1 U1419 ( .A(g369), .Y(n1051) );
  INVX1 U1420 ( .A(g1218), .Y(n1129) );
  INVX1 U1421 ( .A(g1400), .Y(n1085) );
  INVX1 U1422 ( .A(g1397), .Y(n1080) );
  INVX1 U1423 ( .A(g758), .Y(n1070) );
  INVX1 U1424 ( .A(g1386), .Y(n1138) );
  INVX1 U1425 ( .A(g207), .Y(n1046) );
  INVX1 U1426 ( .A(g213), .Y(n1119) );
  INVX1 U1427 ( .A(g186), .Y(n1068) );
  INVX1 U1428 ( .A(g1377), .Y(n1118) );
  INVX1 U1429 ( .A(g1383), .Y(n1087) );
  INVX1 U1430 ( .A(g1371), .Y(n1061) );
  INVX1 U1431 ( .A(g1365), .Y(n1077) );
  INVX1 U1432 ( .A(g1380), .Y(n1154) );
  INVX1 U1433 ( .A(g865), .Y(n1101) );
  INVX1 U1434 ( .A(g877), .Y(n1317) );
  INVX1 U1435 ( .A(g82), .Y(n1384) );
  INVX1 U1436 ( .A(g1810), .Y(g5816) );
  INVX1 U1437 ( .A(g23), .Y(g3327) );
endmodule

